-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 12 2017 08:26:01

-- File Generated:     Dec 6 2018 15:12:25

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "uart" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of uart
entity uart is
port (
    output_axis_tdata : out std_logic_vector(7 downto 0);
    input_axis_tdata : in std_logic_vector(7 downto 0);
    txd : out std_logic;
    tx_busy : out std_logic;
    rxd : in std_logic;
    rx_overrun_error : out std_logic;
    rx_frame_error : out std_logic;
    rx_busy : out std_logic;
    rst : in std_logic;
    output_axis_tvalid : out std_logic;
    output_axis_tready : in std_logic;
    input_axis_tvalid : in std_logic;
    input_axis_tready : out std_logic;
    clk : in std_logic);
end uart;

-- Architecture of uart
-- View name is \INTERFACE\
architecture \INTERFACE\ of uart is

signal \N__9136\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9114\ : std_logic;
signal \N__9107\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9088\ : std_logic;
signal \N__9087\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9078\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9061\ : std_logic;
signal \N__9060\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9051\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9043\ : std_logic;
signal \N__9042\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9033\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9024\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8989\ : std_logic;
signal \N__8988\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8980\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8971\ : std_logic;
signal \N__8970\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8962\ : std_logic;
signal \N__8961\ : std_logic;
signal \N__8954\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8944\ : std_logic;
signal \N__8943\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8934\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8926\ : std_logic;
signal \N__8925\ : std_logic;
signal \N__8918\ : std_logic;
signal \N__8917\ : std_logic;
signal \N__8916\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8907\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8898\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8889\ : std_logic;
signal \N__8872\ : std_logic;
signal \N__8871\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8859\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8852\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8848\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8839\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8835\ : std_logic;
signal \N__8832\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8824\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8803\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8799\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8793\ : std_logic;
signal \N__8790\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8782\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8775\ : std_logic;
signal \N__8772\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8757\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8748\ : std_logic;
signal \N__8745\ : std_logic;
signal \N__8742\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8738\ : std_logic;
signal \N__8735\ : std_logic;
signal \N__8730\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8724\ : std_logic;
signal \N__8721\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8713\ : std_logic;
signal \N__8710\ : std_logic;
signal \N__8701\ : std_logic;
signal \N__8698\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8694\ : std_logic;
signal \N__8691\ : std_logic;
signal \N__8688\ : std_logic;
signal \N__8685\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8674\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8668\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8626\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8604\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8595\ : std_logic;
signal \N__8592\ : std_logic;
signal \N__8589\ : std_logic;
signal \N__8586\ : std_logic;
signal \N__8583\ : std_logic;
signal \N__8578\ : std_logic;
signal \N__8575\ : std_logic;
signal \N__8572\ : std_logic;
signal \N__8571\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8566\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8558\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8532\ : std_logic;
signal \N__8529\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8515\ : std_logic;
signal \N__8512\ : std_logic;
signal \N__8509\ : std_logic;
signal \N__8506\ : std_logic;
signal \N__8503\ : std_logic;
signal \N__8500\ : std_logic;
signal \N__8491\ : std_logic;
signal \N__8488\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8484\ : std_logic;
signal \N__8481\ : std_logic;
signal \N__8478\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8470\ : std_logic;
signal \N__8467\ : std_logic;
signal \N__8464\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8458\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8454\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8434\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8382\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8379\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8376\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8367\ : std_logic;
signal \N__8366\ : std_logic;
signal \N__8363\ : std_logic;
signal \N__8360\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8356\ : std_logic;
signal \N__8355\ : std_logic;
signal \N__8352\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8348\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8344\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8335\ : std_logic;
signal \N__8334\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8332\ : std_logic;
signal \N__8331\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8329\ : std_logic;
signal \N__8328\ : std_logic;
signal \N__8315\ : std_logic;
signal \N__8298\ : std_logic;
signal \N__8291\ : std_logic;
signal \N__8288\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8270\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8268\ : std_logic;
signal \N__8267\ : std_logic;
signal \N__8266\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8264\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8262\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8259\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8256\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8248\ : std_logic;
signal \N__8247\ : std_logic;
signal \N__8246\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8244\ : std_logic;
signal \N__8243\ : std_logic;
signal \N__8242\ : std_logic;
signal \N__8241\ : std_logic;
signal \N__8238\ : std_logic;
signal \N__8233\ : std_logic;
signal \N__8224\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8208\ : std_logic;
signal \N__8199\ : std_logic;
signal \N__8196\ : std_logic;
signal \N__8189\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8175\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8169\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8150\ : std_logic;
signal \N__8147\ : std_logic;
signal \N__8144\ : std_logic;
signal \N__8141\ : std_logic;
signal \N__8134\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8130\ : std_logic;
signal \N__8127\ : std_logic;
signal \N__8124\ : std_logic;
signal \N__8121\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8110\ : std_logic;
signal \N__8107\ : std_logic;
signal \N__8106\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8097\ : std_logic;
signal \N__8094\ : std_logic;
signal \N__8091\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8083\ : std_logic;
signal \N__8080\ : std_logic;
signal \N__8079\ : std_logic;
signal \N__8076\ : std_logic;
signal \N__8073\ : std_logic;
signal \N__8070\ : std_logic;
signal \N__8067\ : std_logic;
signal \N__8062\ : std_logic;
signal \N__8059\ : std_logic;
signal \N__8056\ : std_logic;
signal \N__8055\ : std_logic;
signal \N__8052\ : std_logic;
signal \N__8049\ : std_logic;
signal \N__8046\ : std_logic;
signal \N__8043\ : std_logic;
signal \N__8040\ : std_logic;
signal \N__8037\ : std_logic;
signal \N__8032\ : std_logic;
signal \N__8029\ : std_logic;
signal \N__8028\ : std_logic;
signal \N__8025\ : std_logic;
signal \N__8022\ : std_logic;
signal \N__8019\ : std_logic;
signal \N__8016\ : std_logic;
signal \N__8013\ : std_logic;
signal \N__8010\ : std_logic;
signal \N__8005\ : std_logic;
signal \N__8002\ : std_logic;
signal \N__7999\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7995\ : std_logic;
signal \N__7992\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7980\ : std_logic;
signal \N__7975\ : std_logic;
signal \N__7972\ : std_logic;
signal \N__7971\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7969\ : std_logic;
signal \N__7966\ : std_logic;
signal \N__7963\ : std_logic;
signal \N__7960\ : std_logic;
signal \N__7959\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7949\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7940\ : std_logic;
signal \N__7939\ : std_logic;
signal \N__7936\ : std_logic;
signal \N__7925\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7917\ : std_logic;
signal \N__7914\ : std_logic;
signal \N__7909\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7905\ : std_logic;
signal \N__7902\ : std_logic;
signal \N__7899\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7891\ : std_logic;
signal \N__7888\ : std_logic;
signal \N__7885\ : std_logic;
signal \N__7884\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7882\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7878\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7874\ : std_logic;
signal \N__7871\ : std_logic;
signal \N__7868\ : std_logic;
signal \N__7865\ : std_logic;
signal \N__7862\ : std_logic;
signal \N__7859\ : std_logic;
signal \N__7856\ : std_logic;
signal \N__7853\ : std_logic;
signal \N__7850\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7846\ : std_logic;
signal \N__7843\ : std_logic;
signal \N__7838\ : std_logic;
signal \N__7831\ : std_logic;
signal \N__7828\ : std_logic;
signal \N__7821\ : std_logic;
signal \N__7818\ : std_logic;
signal \N__7813\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7806\ : std_logic;
signal \N__7803\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7792\ : std_logic;
signal \N__7789\ : std_logic;
signal \N__7788\ : std_logic;
signal \N__7787\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7785\ : std_logic;
signal \N__7784\ : std_logic;
signal \N__7781\ : std_logic;
signal \N__7778\ : std_logic;
signal \N__7775\ : std_logic;
signal \N__7772\ : std_logic;
signal \N__7769\ : std_logic;
signal \N__7766\ : std_logic;
signal \N__7763\ : std_logic;
signal \N__7760\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7750\ : std_logic;
signal \N__7747\ : std_logic;
signal \N__7744\ : std_logic;
signal \N__7735\ : std_logic;
signal \N__7732\ : std_logic;
signal \N__7729\ : std_logic;
signal \N__7724\ : std_logic;
signal \N__7721\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7711\ : std_logic;
signal \N__7708\ : std_logic;
signal \N__7707\ : std_logic;
signal \N__7704\ : std_logic;
signal \N__7701\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7693\ : std_logic;
signal \N__7690\ : std_logic;
signal \N__7687\ : std_logic;
signal \N__7684\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7675\ : std_logic;
signal \N__7672\ : std_logic;
signal \N__7669\ : std_logic;
signal \N__7666\ : std_logic;
signal \N__7663\ : std_logic;
signal \N__7660\ : std_logic;
signal \N__7659\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7657\ : std_logic;
signal \N__7656\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7654\ : std_logic;
signal \N__7653\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7651\ : std_logic;
signal \N__7650\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7645\ : std_logic;
signal \N__7642\ : std_logic;
signal \N__7639\ : std_logic;
signal \N__7622\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7608\ : std_logic;
signal \N__7607\ : std_logic;
signal \N__7606\ : std_logic;
signal \N__7605\ : std_logic;
signal \N__7602\ : std_logic;
signal \N__7595\ : std_logic;
signal \N__7592\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7575\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7567\ : std_logic;
signal \N__7564\ : std_logic;
signal \N__7563\ : std_logic;
signal \N__7560\ : std_logic;
signal \N__7557\ : std_logic;
signal \N__7552\ : std_logic;
signal \N__7549\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7543\ : std_logic;
signal \N__7540\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7531\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7526\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7524\ : std_logic;
signal \N__7523\ : std_logic;
signal \N__7522\ : std_logic;
signal \N__7521\ : std_logic;
signal \N__7520\ : std_logic;
signal \N__7519\ : std_logic;
signal \N__7518\ : std_logic;
signal \N__7515\ : std_logic;
signal \N__7498\ : std_logic;
signal \N__7493\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7487\ : std_logic;
signal \N__7486\ : std_logic;
signal \N__7485\ : std_logic;
signal \N__7484\ : std_logic;
signal \N__7483\ : std_logic;
signal \N__7482\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7478\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7456\ : std_logic;
signal \N__7441\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7437\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7433\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7431\ : std_logic;
signal \N__7430\ : std_logic;
signal \N__7425\ : std_logic;
signal \N__7422\ : std_logic;
signal \N__7419\ : std_logic;
signal \N__7414\ : std_logic;
signal \N__7405\ : std_logic;
signal \N__7402\ : std_logic;
signal \N__7399\ : std_logic;
signal \N__7396\ : std_logic;
signal \N__7393\ : std_logic;
signal \N__7390\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7382\ : std_logic;
signal \N__7381\ : std_logic;
signal \N__7380\ : std_logic;
signal \N__7379\ : std_logic;
signal \N__7378\ : std_logic;
signal \N__7377\ : std_logic;
signal \N__7376\ : std_logic;
signal \N__7375\ : std_logic;
signal \N__7374\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7372\ : std_logic;
signal \N__7371\ : std_logic;
signal \N__7370\ : std_logic;
signal \N__7369\ : std_logic;
signal \N__7368\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7366\ : std_logic;
signal \N__7365\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7362\ : std_logic;
signal \N__7361\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7359\ : std_logic;
signal \N__7358\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7356\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7353\ : std_logic;
signal \N__7352\ : std_logic;
signal \N__7285\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7279\ : std_logic;
signal \N__7276\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7270\ : std_logic;
signal \N__7267\ : std_logic;
signal \N__7266\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7263\ : std_logic;
signal \N__7262\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7256\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7254\ : std_logic;
signal \N__7253\ : std_logic;
signal \N__7252\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7245\ : std_logic;
signal \N__7244\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7242\ : std_logic;
signal \N__7241\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7239\ : std_logic;
signal \N__7238\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7236\ : std_logic;
signal \N__7233\ : std_logic;
signal \N__7232\ : std_logic;
signal \N__7231\ : std_logic;
signal \N__7228\ : std_logic;
signal \N__7227\ : std_logic;
signal \N__7224\ : std_logic;
signal \N__7221\ : std_logic;
signal \N__7218\ : std_logic;
signal \N__7215\ : std_logic;
signal \N__7212\ : std_logic;
signal \N__7209\ : std_logic;
signal \N__7206\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7200\ : std_logic;
signal \N__7197\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7188\ : std_logic;
signal \N__7187\ : std_logic;
signal \N__7186\ : std_logic;
signal \N__7185\ : std_logic;
signal \N__7182\ : std_logic;
signal \N__7181\ : std_logic;
signal \N__7178\ : std_logic;
signal \N__7177\ : std_logic;
signal \N__7176\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7172\ : std_logic;
signal \N__7169\ : std_logic;
signal \N__7164\ : std_logic;
signal \N__7163\ : std_logic;
signal \N__7162\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7158\ : std_logic;
signal \N__7155\ : std_logic;
signal \N__7152\ : std_logic;
signal \N__7149\ : std_logic;
signal \N__7140\ : std_logic;
signal \N__7137\ : std_logic;
signal \N__7134\ : std_logic;
signal \N__7133\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7118\ : std_logic;
signal \N__7115\ : std_logic;
signal \N__7108\ : std_logic;
signal \N__7105\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7096\ : std_logic;
signal \N__7093\ : std_logic;
signal \N__7090\ : std_logic;
signal \N__7087\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7074\ : std_logic;
signal \N__7073\ : std_logic;
signal \N__7072\ : std_logic;
signal \N__7069\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7061\ : std_logic;
signal \N__7054\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7037\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7023\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7008\ : std_logic;
signal \N__7005\ : std_logic;
signal \N__7002\ : std_logic;
signal \N__6999\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6981\ : std_logic;
signal \N__6974\ : std_logic;
signal \N__6961\ : std_logic;
signal \N__6960\ : std_logic;
signal \N__6957\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6951\ : std_logic;
signal \N__6948\ : std_logic;
signal \N__6945\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6930\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6924\ : std_logic;
signal \N__6921\ : std_logic;
signal \N__6918\ : std_logic;
signal \N__6915\ : std_logic;
signal \N__6912\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6904\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6898\ : std_logic;
signal \N__6897\ : std_logic;
signal \N__6894\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6877\ : std_logic;
signal \N__6874\ : std_logic;
signal \N__6873\ : std_logic;
signal \N__6870\ : std_logic;
signal \N__6867\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6856\ : std_logic;
signal \N__6853\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6849\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6838\ : std_logic;
signal \N__6837\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6834\ : std_logic;
signal \N__6833\ : std_logic;
signal \N__6832\ : std_logic;
signal \N__6827\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6821\ : std_logic;
signal \N__6816\ : std_logic;
signal \N__6813\ : std_logic;
signal \N__6812\ : std_logic;
signal \N__6811\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6809\ : std_logic;
signal \N__6808\ : std_logic;
signal \N__6807\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6805\ : std_logic;
signal \N__6804\ : std_logic;
signal \N__6799\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6787\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6777\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6774\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6756\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6733\ : std_logic;
signal \N__6730\ : std_logic;
signal \N__6727\ : std_logic;
signal \N__6726\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6723\ : std_logic;
signal \N__6722\ : std_logic;
signal \N__6721\ : std_logic;
signal \N__6714\ : std_logic;
signal \N__6713\ : std_logic;
signal \N__6712\ : std_logic;
signal \N__6711\ : std_logic;
signal \N__6710\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6708\ : std_logic;
signal \N__6707\ : std_logic;
signal \N__6700\ : std_logic;
signal \N__6699\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6696\ : std_logic;
signal \N__6693\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6691\ : std_logic;
signal \N__6690\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6677\ : std_logic;
signal \N__6670\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6668\ : std_logic;
signal \N__6667\ : std_logic;
signal \N__6664\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6643\ : std_logic;
signal \N__6638\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6632\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6603\ : std_logic;
signal \N__6598\ : std_logic;
signal \N__6597\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6594\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6574\ : std_logic;
signal \N__6573\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6570\ : std_logic;
signal \N__6569\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6567\ : std_logic;
signal \N__6566\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6560\ : std_logic;
signal \N__6555\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6539\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6533\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6495\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6477\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6466\ : std_logic;
signal \N__6465\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6461\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6451\ : std_logic;
signal \N__6448\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6431\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6421\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6412\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6406\ : std_logic;
signal \N__6403\ : std_logic;
signal \N__6400\ : std_logic;
signal \N__6397\ : std_logic;
signal \N__6394\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6388\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6382\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6370\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6349\ : std_logic;
signal \N__6346\ : std_logic;
signal \N__6343\ : std_logic;
signal \N__6340\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6325\ : std_logic;
signal \N__6322\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6320\ : std_logic;
signal \N__6315\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6312\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6304\ : std_logic;
signal \N__6303\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6300\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6297\ : std_logic;
signal \N__6296\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6294\ : std_logic;
signal \N__6293\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6288\ : std_logic;
signal \N__6287\ : std_logic;
signal \N__6282\ : std_logic;
signal \N__6279\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6273\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6237\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6208\ : std_logic;
signal \N__6207\ : std_logic;
signal \N__6204\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6193\ : std_logic;
signal \N__6190\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6172\ : std_logic;
signal \N__6169\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6163\ : std_logic;
signal \N__6160\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6154\ : std_logic;
signal \N__6151\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6145\ : std_logic;
signal \N__6142\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6124\ : std_logic;
signal \N__6121\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6109\ : std_logic;
signal \N__6106\ : std_logic;
signal \N__6103\ : std_logic;
signal \N__6100\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6091\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6063\ : std_logic;
signal \N__6060\ : std_logic;
signal \N__6057\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6027\ : std_logic;
signal \N__6024\ : std_logic;
signal \N__6021\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5997\ : std_logic;
signal \N__5994\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5985\ : std_logic;
signal \N__5982\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5962\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5929\ : std_logic;
signal \N__5928\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5922\ : std_logic;
signal \N__5919\ : std_logic;
signal \N__5916\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5910\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5896\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5881\ : std_logic;
signal \N__5878\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5869\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5854\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5844\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5836\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5820\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5809\ : std_logic;
signal \N__5806\ : std_logic;
signal \N__5803\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5791\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5754\ : std_logic;
signal \N__5751\ : std_logic;
signal \N__5748\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5721\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5715\ : std_logic;
signal \N__5712\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5704\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5695\ : std_logic;
signal \N__5692\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5685\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5674\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5658\ : std_logic;
signal \N__5655\ : std_logic;
signal \N__5652\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5622\ : std_logic;
signal \N__5619\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5610\ : std_logic;
signal \N__5607\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5586\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5577\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5554\ : std_logic;
signal \N__5553\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5539\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5526\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5519\ : std_logic;
signal \N__5516\ : std_logic;
signal \N__5511\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5464\ : std_logic;
signal \N__5461\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5454\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5431\ : std_logic;
signal \N__5428\ : std_logic;
signal \N__5425\ : std_logic;
signal \N__5422\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5418\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5412\ : std_logic;
signal \N__5409\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5390\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5374\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5364\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5361\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5355\ : std_logic;
signal \N__5348\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5320\ : std_logic;
signal \N__5317\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5296\ : std_logic;
signal \N__5295\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5286\ : std_logic;
signal \N__5283\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5269\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5230\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5218\ : std_logic;
signal \N__5215\ : std_logic;
signal \N__5212\ : std_logic;
signal \N__5209\ : std_logic;
signal \N__5206\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5173\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5163\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5150\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5128\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5108\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5095\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5086\ : std_logic;
signal \N__5083\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5071\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5053\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5035\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5026\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5020\ : std_logic;
signal \N__5017\ : std_logic;
signal \N__5014\ : std_logic;
signal \N__5013\ : std_logic;
signal \N__5010\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__4999\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4993\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4978\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4969\ : std_logic;
signal \N__4966\ : std_logic;
signal \N__4963\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4951\ : std_logic;
signal \N__4948\ : std_logic;
signal \N__4945\ : std_logic;
signal \N__4942\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4940\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4936\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4933\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4921\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4913\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4906\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4874\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4852\ : std_logic;
signal \N__4849\ : std_logic;
signal \N__4848\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4842\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4816\ : std_logic;
signal \N__4813\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4804\ : std_logic;
signal \N__4801\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4795\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4768\ : std_logic;
signal \N__4765\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4759\ : std_logic;
signal \N__4758\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4707\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4683\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4675\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4668\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4641\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4621\ : std_logic;
signal \N__4618\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4606\ : std_logic;
signal \N__4603\ : std_logic;
signal \N__4600\ : std_logic;
signal \N__4597\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4594\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4576\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4552\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4540\ : std_logic;
signal \N__4537\ : std_logic;
signal \N__4534\ : std_logic;
signal \N__4531\ : std_logic;
signal \N__4528\ : std_logic;
signal \N__4525\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4518\ : std_logic;
signal \N__4515\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4495\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4488\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4474\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4455\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4447\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4423\ : std_logic;
signal \N__4420\ : std_logic;
signal \N__4417\ : std_logic;
signal \N__4414\ : std_logic;
signal \N__4411\ : std_logic;
signal \N__4408\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4399\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4395\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4384\ : std_logic;
signal \N__4381\ : std_logic;
signal \N__4378\ : std_logic;
signal \N__4375\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4369\ : std_logic;
signal \N__4368\ : std_logic;
signal \N__4365\ : std_logic;
signal \N__4362\ : std_logic;
signal \N__4357\ : std_logic;
signal \N__4354\ : std_logic;
signal \N__4351\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4347\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4321\ : std_logic;
signal \N__4318\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4306\ : std_logic;
signal \N__4303\ : std_logic;
signal \N__4300\ : std_logic;
signal \N__4297\ : std_logic;
signal \N__4294\ : std_logic;
signal \N__4291\ : std_logic;
signal \N__4288\ : std_logic;
signal \N__4285\ : std_logic;
signal \N__4282\ : std_logic;
signal \N__4279\ : std_logic;
signal \N__4276\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4270\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4264\ : std_logic;
signal \N__4263\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4261\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4239\ : std_logic;
signal \N__4236\ : std_logic;
signal \N__4229\ : std_logic;
signal \N__4226\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4212\ : std_logic;
signal \N__4211\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4207\ : std_logic;
signal \N__4206\ : std_logic;
signal \N__4201\ : std_logic;
signal \N__4198\ : std_logic;
signal \N__4195\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4189\ : std_logic;
signal \N__4180\ : std_logic;
signal \N__4177\ : std_logic;
signal \N__4174\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4170\ : std_logic;
signal \N__4167\ : std_logic;
signal \N__4162\ : std_logic;
signal \N__4161\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4159\ : std_logic;
signal \N__4156\ : std_logic;
signal \N__4149\ : std_logic;
signal \N__4144\ : std_logic;
signal \N__4141\ : std_logic;
signal \N__4138\ : std_logic;
signal \N__4135\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4131\ : std_logic;
signal \N__4128\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4120\ : std_logic;
signal \N__4117\ : std_logic;
signal \N__4114\ : std_logic;
signal \N__4111\ : std_logic;
signal \N__4104\ : std_logic;
signal \N__4099\ : std_logic;
signal \N__4098\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4092\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4086\ : std_logic;
signal \N__4083\ : std_logic;
signal \N__4080\ : std_logic;
signal \N__4075\ : std_logic;
signal \N__4074\ : std_logic;
signal \N__4071\ : std_logic;
signal \N__4068\ : std_logic;
signal \N__4065\ : std_logic;
signal \N__4062\ : std_logic;
signal \N__4057\ : std_logic;
signal \N__4054\ : std_logic;
signal \N__4051\ : std_logic;
signal \N__4048\ : std_logic;
signal \N__4045\ : std_logic;
signal \N__4042\ : std_logic;
signal \N__4039\ : std_logic;
signal \N__4036\ : std_logic;
signal \N__4033\ : std_logic;
signal \N__4030\ : std_logic;
signal \N__4029\ : std_logic;
signal \N__4028\ : std_logic;
signal \N__4027\ : std_logic;
signal \N__4024\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4013\ : std_logic;
signal \N__4006\ : std_logic;
signal \N__4003\ : std_logic;
signal \N__4000\ : std_logic;
signal \N__3999\ : std_logic;
signal \N__3998\ : std_logic;
signal \N__3997\ : std_logic;
signal \N__3994\ : std_logic;
signal \N__3989\ : std_logic;
signal \N__3986\ : std_logic;
signal \N__3979\ : std_logic;
signal \N__3976\ : std_logic;
signal \N__3973\ : std_logic;
signal \N__3972\ : std_logic;
signal \N__3969\ : std_logic;
signal \N__3966\ : std_logic;
signal \N__3961\ : std_logic;
signal \N__3960\ : std_logic;
signal \N__3957\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3949\ : std_logic;
signal \N__3946\ : std_logic;
signal \N__3943\ : std_logic;
signal \N__3942\ : std_logic;
signal \N__3939\ : std_logic;
signal \N__3936\ : std_logic;
signal \N__3931\ : std_logic;
signal \N__3930\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3926\ : std_logic;
signal \N__3925\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3923\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3917\ : std_logic;
signal \N__3912\ : std_logic;
signal \N__3909\ : std_logic;
signal \N__3906\ : std_logic;
signal \N__3895\ : std_logic;
signal \N__3894\ : std_logic;
signal \N__3893\ : std_logic;
signal \N__3892\ : std_logic;
signal \N__3891\ : std_logic;
signal \N__3888\ : std_logic;
signal \N__3885\ : std_logic;
signal \N__3880\ : std_logic;
signal \N__3877\ : std_logic;
signal \N__3868\ : std_logic;
signal \N__3867\ : std_logic;
signal \N__3864\ : std_logic;
signal \N__3861\ : std_logic;
signal \N__3858\ : std_logic;
signal \N__3855\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3851\ : std_logic;
signal \N__3848\ : std_logic;
signal \N__3845\ : std_logic;
signal \N__3838\ : std_logic;
signal \N__3835\ : std_logic;
signal \N__3832\ : std_logic;
signal \N__3829\ : std_logic;
signal \N__3826\ : std_logic;
signal \N__3823\ : std_logic;
signal \N__3822\ : std_logic;
signal \N__3821\ : std_logic;
signal \N__3820\ : std_logic;
signal \N__3819\ : std_logic;
signal \N__3818\ : std_logic;
signal \N__3817\ : std_logic;
signal \N__3816\ : std_logic;
signal \N__3815\ : std_logic;
signal \N__3814\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3812\ : std_logic;
signal \N__3811\ : std_logic;
signal \N__3810\ : std_logic;
signal \N__3809\ : std_logic;
signal \N__3808\ : std_logic;
signal \N__3807\ : std_logic;
signal \N__3806\ : std_logic;
signal \N__3805\ : std_logic;
signal \N__3804\ : std_logic;
signal \N__3803\ : std_logic;
signal \N__3800\ : std_logic;
signal \N__3799\ : std_logic;
signal \N__3796\ : std_logic;
signal \N__3779\ : std_logic;
signal \N__3766\ : std_logic;
signal \N__3761\ : std_logic;
signal \N__3750\ : std_logic;
signal \N__3739\ : std_logic;
signal \N__3738\ : std_logic;
signal \N__3735\ : std_logic;
signal \N__3734\ : std_logic;
signal \N__3733\ : std_logic;
signal \N__3730\ : std_logic;
signal \N__3727\ : std_logic;
signal \N__3724\ : std_logic;
signal \N__3721\ : std_logic;
signal \N__3712\ : std_logic;
signal \N__3709\ : std_logic;
signal \N__3706\ : std_logic;
signal \N__3703\ : std_logic;
signal \N__3700\ : std_logic;
signal \N__3697\ : std_logic;
signal \N__3696\ : std_logic;
signal \N__3695\ : std_logic;
signal \N__3694\ : std_logic;
signal \N__3691\ : std_logic;
signal \N__3690\ : std_logic;
signal \N__3689\ : std_logic;
signal \N__3686\ : std_logic;
signal \N__3683\ : std_logic;
signal \N__3682\ : std_logic;
signal \N__3675\ : std_logic;
signal \N__3666\ : std_logic;
signal \N__3661\ : std_logic;
signal \N__3660\ : std_logic;
signal \N__3659\ : std_logic;
signal \N__3658\ : std_logic;
signal \N__3657\ : std_logic;
signal \N__3656\ : std_logic;
signal \N__3649\ : std_logic;
signal \N__3642\ : std_logic;
signal \N__3637\ : std_logic;
signal \N__3634\ : std_logic;
signal \N__3631\ : std_logic;
signal \N__3628\ : std_logic;
signal \N__3625\ : std_logic;
signal \N__3622\ : std_logic;
signal \N__3619\ : std_logic;
signal \N__3616\ : std_logic;
signal \N__3613\ : std_logic;
signal \N__3610\ : std_logic;
signal \N__3607\ : std_logic;
signal \N__3604\ : std_logic;
signal \N__3601\ : std_logic;
signal \N__3600\ : std_logic;
signal \N__3599\ : std_logic;
signal \N__3596\ : std_logic;
signal \N__3593\ : std_logic;
signal \N__3590\ : std_logic;
signal \N__3583\ : std_logic;
signal \N__3582\ : std_logic;
signal \N__3579\ : std_logic;
signal \N__3576\ : std_logic;
signal \N__3573\ : std_logic;
signal \N__3568\ : std_logic;
signal \N__3565\ : std_logic;
signal \N__3562\ : std_logic;
signal \N__3559\ : std_logic;
signal \N__3556\ : std_logic;
signal \N__3555\ : std_logic;
signal \N__3552\ : std_logic;
signal \N__3551\ : std_logic;
signal \N__3550\ : std_logic;
signal \N__3549\ : std_logic;
signal \N__3548\ : std_logic;
signal \N__3545\ : std_logic;
signal \N__3542\ : std_logic;
signal \N__3539\ : std_logic;
signal \N__3536\ : std_logic;
signal \N__3533\ : std_logic;
signal \N__3528\ : std_logic;
signal \N__3517\ : std_logic;
signal \N__3514\ : std_logic;
signal \N__3511\ : std_logic;
signal \N__3508\ : std_logic;
signal \N__3507\ : std_logic;
signal \N__3506\ : std_logic;
signal \N__3505\ : std_logic;
signal \N__3504\ : std_logic;
signal \N__3503\ : std_logic;
signal \N__3502\ : std_logic;
signal \N__3499\ : std_logic;
signal \N__3494\ : std_logic;
signal \N__3485\ : std_logic;
signal \N__3478\ : std_logic;
signal \N__3475\ : std_logic;
signal \N__3472\ : std_logic;
signal \N__3469\ : std_logic;
signal \N__3466\ : std_logic;
signal \N__3463\ : std_logic;
signal \N__3460\ : std_logic;
signal \N__3457\ : std_logic;
signal \N__3454\ : std_logic;
signal \N__3451\ : std_logic;
signal \N__3448\ : std_logic;
signal \N__3445\ : std_logic;
signal \N__3442\ : std_logic;
signal \N__3439\ : std_logic;
signal \N__3436\ : std_logic;
signal \N__3435\ : std_logic;
signal \N__3432\ : std_logic;
signal \N__3429\ : std_logic;
signal \N__3424\ : std_logic;
signal \N__3421\ : std_logic;
signal \N__3418\ : std_logic;
signal \N__3415\ : std_logic;
signal \N__3412\ : std_logic;
signal \N__3409\ : std_logic;
signal \N__3406\ : std_logic;
signal \N__3405\ : std_logic;
signal \N__3402\ : std_logic;
signal \N__3399\ : std_logic;
signal \N__3394\ : std_logic;
signal \N__3393\ : std_logic;
signal \N__3390\ : std_logic;
signal \N__3387\ : std_logic;
signal \N__3382\ : std_logic;
signal \N__3379\ : std_logic;
signal \N__3376\ : std_logic;
signal \N__3373\ : std_logic;
signal \N__3370\ : std_logic;
signal \N__3367\ : std_logic;
signal \N__3364\ : std_logic;
signal \N__3361\ : std_logic;
signal \N__3358\ : std_logic;
signal \N__3355\ : std_logic;
signal \N__3352\ : std_logic;
signal \N__3351\ : std_logic;
signal \N__3348\ : std_logic;
signal \N__3345\ : std_logic;
signal \N__3340\ : std_logic;
signal \N__3337\ : std_logic;
signal \N__3334\ : std_logic;
signal \N__3331\ : std_logic;
signal \N__3328\ : std_logic;
signal \N__3325\ : std_logic;
signal \N__3322\ : std_logic;
signal \N__3319\ : std_logic;
signal \N__3316\ : std_logic;
signal \N__3313\ : std_logic;
signal \N__3310\ : std_logic;
signal \N__3307\ : std_logic;
signal \N__3304\ : std_logic;
signal \N__3301\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal tx_busy_c : std_logic;
signal \uart_tx_inst.n721\ : std_logic;
signal input_axis_tready_c : std_logic;
signal \uart_tx_inst.n701\ : std_logic;
signal \uart_tx_inst.n535\ : std_logic;
signal rx_busy_c : std_logic;
signal \n588_cascade_\ : std_logic;
signal \n707_cascade_\ : std_logic;
signal \uart_tx_inst.n7_cascade_\ : std_logic;
signal n1165 : std_logic;
signal n4 : std_logic;
signal \uart_tx_inst.n613\ : std_logic;
signal n707 : std_logic;
signal rx_overrun_error_c : std_logic;
signal \uart_rx_inst.n984\ : std_logic;
signal \n705_cascade_\ : std_logic;
signal \n1167_cascade_\ : std_logic;
signal n1698 : std_logic;
signal \uart_rx_inst.n677_cascade_\ : std_logic;
signal \uart_rx_inst.n607_cascade_\ : std_logic;
signal \uart_rx_inst.n603_cascade_\ : std_logic;
signal n1471 : std_logic;
signal \uart_tx_inst.n485_cascade_\ : std_logic;
signal \uart_tx_inst.n30_adj_196_cascade_\ : std_logic;
signal \uart_tx_inst.n34_cascade_\ : std_logic;
signal \uart_tx_inst.n189_cascade_\ : std_logic;
signal \uart_tx_inst.bit_cnt_0\ : std_logic;
signal \uart_tx_inst.n7_adj_195\ : std_logic;
signal \uart_tx_inst.bit_cnt_1\ : std_logic;
signal \uart_tx_inst.n15_cascade_\ : std_logic;
signal bit_cnt_2 : std_logic;
signal \uart_tx_inst.bit_cnt_3\ : std_logic;
signal \uart_tx_inst.n1723_cascade_\ : std_logic;
signal \uart_rx_inst.n681\ : std_logic;
signal \uart_tx_inst.n13\ : std_logic;
signal output_axis_tready_c : std_logic;
signal output_axis_tvalid_c : std_logic;
signal \uart_rx_inst.n30_cascade_\ : std_logic;
signal \uart_rx_inst.n32_cascade_\ : std_logic;
signal \uart_rx_inst.n34\ : std_logic;
signal \output_axis_tvalid_N_175_cascade_\ : std_logic;
signal \uart_rx_inst.n509_cascade_\ : std_logic;
signal \uart_rx_inst.n31\ : std_logic;
signal \uart_rx_inst.n33\ : std_logic;
signal \uart_rx_inst.n1479\ : std_logic;
signal \uart_rx_inst.n1045\ : std_logic;
signal \uart_rx_inst.output_axis_tvalid_N_174\ : std_logic;
signal \n1711_cascade_\ : std_logic;
signal \n1220_cascade_\ : std_logic;
signal \uart_rx_inst.bit_cnt_3\ : std_logic;
signal \uart_rx_inst.output_axis_tvalid_N_172_cascade_\ : std_logic;
signal \uart_rx_inst.n232_cascade_\ : std_logic;
signal \uart_rx_inst.n1468\ : std_logic;
signal \uart_rx_inst.n1502\ : std_logic;
signal \uart_rx_inst.n235\ : std_logic;
signal \uart_rx_inst.bit_cnt_1\ : std_logic;
signal \uart_rx_inst.bit_cnt_2\ : std_logic;
signal n705 : std_logic;
signal n1167 : std_logic;
signal bit_cnt_0 : std_logic;
signal \uart_rx_inst.n677\ : std_logic;
signal \uart_rx_inst.output_axis_tvalid_N_172\ : std_logic;
signal \uart_rx_inst.output_axis_tvalid_N_173\ : std_logic;
signal \n695_cascade_\ : std_logic;
signal n695 : std_logic;
signal \output_axis_tvalid_N_175\ : std_logic;
signal n680 : std_logic;
signal data_reg_0 : std_logic;
signal output_axis_tdata_c_0 : std_logic;
signal rxd_c : std_logic;
signal \uart_tx_inst.n910_cascade_\ : std_logic;
signal \uart_tx_inst.n920_cascade_\ : std_logic;
signal \uart_tx_inst.n930_cascade_\ : std_logic;
signal \uart_tx_inst.n31_adj_199\ : std_logic;
signal \uart_tx_inst.n915\ : std_logic;
signal \uart_tx_inst.n875_cascade_\ : std_logic;
signal \uart_tx_inst.n880_cascade_\ : std_logic;
signal \uart_tx_inst.n895_cascade_\ : std_logic;
signal \uart_tx_inst.n900_cascade_\ : std_logic;
signal \uart_tx_inst.n925\ : std_logic;
signal \uart_tx_inst.n935\ : std_logic;
signal \uart_rx_inst.n509\ : std_logic;
signal \uart_rx_inst.prescale_reg_0\ : std_logic;
signal \bfn_9_5_0_\ : std_logic;
signal \uart_rx_inst.n1648\ : std_logic;
signal \uart_rx_inst.n1141\ : std_logic;
signal \uart_rx_inst.prescale_reg_1\ : std_logic;
signal \uart_rx_inst.n819\ : std_logic;
signal \uart_rx_inst.n1564\ : std_logic;
signal \uart_rx_inst.prescale_reg_2\ : std_logic;
signal \uart_rx_inst.n814\ : std_logic;
signal \uart_rx_inst.n1565\ : std_logic;
signal \uart_rx_inst.prescale_reg_3\ : std_logic;
signal \uart_rx_inst.n809\ : std_logic;
signal \uart_rx_inst.n1566\ : std_logic;
signal \uart_rx_inst.prescale_reg_4\ : std_logic;
signal \uart_rx_inst.n804\ : std_logic;
signal \uart_rx_inst.n1567\ : std_logic;
signal \uart_rx_inst.n1756\ : std_logic;
signal \uart_rx_inst.prescale_reg_5\ : std_logic;
signal \uart_rx_inst.n799\ : std_logic;
signal \uart_rx_inst.n1568\ : std_logic;
signal \uart_rx_inst.prescale_reg_6\ : std_logic;
signal \uart_rx_inst.n794\ : std_logic;
signal \uart_rx_inst.n1569\ : std_logic;
signal \uart_rx_inst.prescale_reg_7\ : std_logic;
signal \uart_rx_inst.n789\ : std_logic;
signal \uart_rx_inst.n1570\ : std_logic;
signal \uart_rx_inst.n1571\ : std_logic;
signal \uart_rx_inst.prescale_reg_8\ : std_logic;
signal \uart_rx_inst.n784\ : std_logic;
signal \bfn_9_6_0_\ : std_logic;
signal \uart_rx_inst.prescale_reg_9\ : std_logic;
signal \uart_rx_inst.n779\ : std_logic;
signal \uart_rx_inst.n1572\ : std_logic;
signal \uart_rx_inst.n1744\ : std_logic;
signal \uart_rx_inst.prescale_reg_10\ : std_logic;
signal \uart_rx_inst.n774\ : std_logic;
signal \uart_rx_inst.n1573\ : std_logic;
signal \uart_rx_inst.prescale_reg_11\ : std_logic;
signal \uart_rx_inst.n769\ : std_logic;
signal \uart_rx_inst.n1574\ : std_logic;
signal \uart_rx_inst.prescale_reg_12\ : std_logic;
signal \uart_rx_inst.n764\ : std_logic;
signal \uart_rx_inst.n1575\ : std_logic;
signal \uart_rx_inst.prescale_reg_13\ : std_logic;
signal \uart_rx_inst.n759\ : std_logic;
signal \uart_rx_inst.n1576\ : std_logic;
signal \uart_rx_inst.prescale_reg_14\ : std_logic;
signal \uart_rx_inst.n754\ : std_logic;
signal \uart_rx_inst.n1577\ : std_logic;
signal \uart_rx_inst.prescale_reg_15\ : std_logic;
signal \uart_rx_inst.n749\ : std_logic;
signal \uart_rx_inst.n1578\ : std_logic;
signal \uart_rx_inst.n1579\ : std_logic;
signal \uart_rx_inst.prescale_reg_16\ : std_logic;
signal \uart_rx_inst.n744\ : std_logic;
signal \bfn_9_7_0_\ : std_logic;
signal \uart_rx_inst.prescale_reg_17\ : std_logic;
signal \uart_rx_inst.n739\ : std_logic;
signal \uart_rx_inst.n1580\ : std_logic;
signal \uart_rx_inst.n712\ : std_logic;
signal \uart_rx_inst.prescale_reg_18\ : std_logic;
signal \uart_rx_inst.n1581\ : std_logic;
signal \uart_rx_inst.n729\ : std_logic;
signal \uart_rx_inst.n1743\ : std_logic;
signal \uart_rx_inst.n1740\ : std_logic;
signal \uart_rx_inst.n1741\ : std_logic;
signal \uart_rx_inst.n1747\ : std_logic;
signal \uart_rx_inst.n1745\ : std_logic;
signal \uart_rx_inst.n1750\ : std_logic;
signal \uart_rx_inst.n1755\ : std_logic;
signal \uart_rx_inst.n1754\ : std_logic;
signal \uart_rx_inst.n1751\ : std_logic;
signal \uart_rx_inst.n1758\ : std_logic;
signal \uart_rx_inst.n1742\ : std_logic;
signal \uart_rx_inst.n1739\ : std_logic;
signal \uart_rx_inst.n1757\ : std_logic;
signal n1711 : std_logic;
signal n1220 : std_logic;
signal rxd_reg : std_logic;
signal rx_frame_error_c : std_logic;
signal n697 : std_logic;
signal data_reg_6 : std_logic;
signal output_axis_tdata_c_6 : std_logic;
signal data_reg_2 : std_logic;
signal output_axis_tdata_c_2 : std_logic;
signal data_reg_7 : std_logic;
signal output_axis_tdata_c_7 : std_logic;
signal data_reg_4 : std_logic;
signal output_axis_tdata_c_4 : std_logic;
signal data_reg_5 : std_logic;
signal output_axis_tdata_c_5 : std_logic;
signal data_reg_1 : std_logic;
signal output_axis_tdata_c_1 : std_logic;
signal data_reg_3 : std_logic;
signal output_axis_tdata_c_3 : std_logic;
signal n703 : std_logic;
signal \uart_tx_inst.n905_cascade_\ : std_logic;
signal \uart_tx_inst.n890_cascade_\ : std_logic;
signal \uart_tx_inst.n33_adj_198\ : std_logic;
signal \uart_tx_inst.n860_cascade_\ : std_logic;
signal \bfn_11_2_0_\ : std_logic;
signal \uart_tx_inst.prescale_reg_1\ : std_logic;
signal \uart_tx_inst.n1546\ : std_logic;
signal \uart_tx_inst.prescale_reg_2\ : std_logic;
signal \uart_tx_inst.n1547\ : std_logic;
signal \uart_tx_inst.n1170\ : std_logic;
signal \uart_tx_inst.prescale_reg_3\ : std_logic;
signal \uart_tx_inst.n33\ : std_logic;
signal \uart_tx_inst.n1548\ : std_logic;
signal \uart_tx_inst.n1549\ : std_logic;
signal \uart_tx_inst.n1550\ : std_logic;
signal \uart_tx_inst.prescale_reg_6\ : std_logic;
signal \uart_tx_inst.n30\ : std_logic;
signal \uart_tx_inst.n1551\ : std_logic;
signal \uart_tx_inst.prescale_reg_7\ : std_logic;
signal \uart_tx_inst.n29\ : std_logic;
signal \uart_tx_inst.n1552\ : std_logic;
signal \uart_tx_inst.n1553\ : std_logic;
signal \bfn_11_3_0_\ : std_logic;
signal \uart_tx_inst.prescale_reg_9\ : std_logic;
signal \uart_tx_inst.n27\ : std_logic;
signal \uart_tx_inst.n1554\ : std_logic;
signal \uart_tx_inst.prescale_reg_10\ : std_logic;
signal \uart_tx_inst.n26\ : std_logic;
signal \uart_tx_inst.n1555\ : std_logic;
signal \uart_tx_inst.prescale_reg_11\ : std_logic;
signal \uart_tx_inst.n25\ : std_logic;
signal \uart_tx_inst.n1556\ : std_logic;
signal \uart_tx_inst.prescale_reg_12\ : std_logic;
signal \uart_tx_inst.n24\ : std_logic;
signal \uart_tx_inst.n1557\ : std_logic;
signal \uart_tx_inst.prescale_reg_13\ : std_logic;
signal \uart_tx_inst.n23\ : std_logic;
signal \uart_tx_inst.n1558\ : std_logic;
signal \uart_tx_inst.prescale_reg_14\ : std_logic;
signal \uart_tx_inst.n22\ : std_logic;
signal \uart_tx_inst.n1559\ : std_logic;
signal \uart_tx_inst.prescale_reg_15\ : std_logic;
signal \uart_tx_inst.n21\ : std_logic;
signal \uart_tx_inst.n1560\ : std_logic;
signal \uart_tx_inst.n1561\ : std_logic;
signal \uart_tx_inst.prescale_reg_16\ : std_logic;
signal \uart_tx_inst.n20\ : std_logic;
signal \bfn_11_4_0_\ : std_logic;
signal \uart_tx_inst.prescale_reg_17\ : std_logic;
signal \uart_tx_inst.n19\ : std_logic;
signal \uart_tx_inst.n1562\ : std_logic;
signal \uart_tx_inst.prescale_reg_18\ : std_logic;
signal \uart_tx_inst.n1563\ : std_logic;
signal \uart_tx_inst.n18\ : std_logic;
signal \uart_rx_inst.n328\ : std_logic;
signal \bfn_11_5_0_\ : std_logic;
signal \uart_rx_inst.n327\ : std_logic;
signal \uart_rx_inst.n1530\ : std_logic;
signal \uart_rx_inst.n326\ : std_logic;
signal \uart_rx_inst.n1531\ : std_logic;
signal \uart_rx_inst.n325\ : std_logic;
signal \uart_rx_inst.n1532\ : std_logic;
signal \uart_rx_inst.n324\ : std_logic;
signal \uart_rx_inst.n1533\ : std_logic;
signal \uart_rx_inst.n323\ : std_logic;
signal \uart_rx_inst.n1534\ : std_logic;
signal \uart_rx_inst.n322\ : std_logic;
signal \uart_rx_inst.n1535\ : std_logic;
signal \uart_rx_inst.n321\ : std_logic;
signal \uart_rx_inst.n1536\ : std_logic;
signal \uart_rx_inst.n1537\ : std_logic;
signal \uart_rx_inst.n320\ : std_logic;
signal \bfn_11_6_0_\ : std_logic;
signal \uart_rx_inst.n319\ : std_logic;
signal \uart_rx_inst.n1538\ : std_logic;
signal \uart_rx_inst.n318\ : std_logic;
signal \uart_rx_inst.n1539\ : std_logic;
signal \uart_rx_inst.n317\ : std_logic;
signal \uart_rx_inst.n1540\ : std_logic;
signal \uart_rx_inst.n316\ : std_logic;
signal \uart_rx_inst.n1541\ : std_logic;
signal \uart_rx_inst.n315\ : std_logic;
signal \uart_rx_inst.n1542\ : std_logic;
signal \uart_rx_inst.n314\ : std_logic;
signal \uart_rx_inst.n1543\ : std_logic;
signal \uart_rx_inst.n313\ : std_logic;
signal \uart_rx_inst.n1544\ : std_logic;
signal \uart_rx_inst.n1545\ : std_logic;
signal \bfn_11_7_0_\ : std_logic;
signal \uart_rx_inst.n312\ : std_logic;
signal \uart_rx_inst.n232\ : std_logic;
signal \uart_rx_inst.n1746\ : std_logic;
signal \uart_tx_inst.prescale_reg_0\ : std_logic;
signal \uart_tx_inst.n32_adj_197\ : std_logic;
signal \uart_tx_inst.n32\ : std_logic;
signal \uart_tx_inst.n865_cascade_\ : std_logic;
signal \uart_tx_inst.prescale_reg_4\ : std_logic;
signal \uart_tx_inst.n31\ : std_logic;
signal \uart_tx_inst.n870_cascade_\ : std_logic;
signal \uart_tx_inst.prescale_reg_5\ : std_logic;
signal \uart_tx_inst.n485\ : std_logic;
signal \uart_tx_inst.n28\ : std_logic;
signal \input_axis_tready_N_72\ : std_logic;
signal \uart_tx_inst.n885_cascade_\ : std_logic;
signal \uart_tx_inst.n165\ : std_logic;
signal \uart_tx_inst.prescale_reg_8\ : std_logic;
signal \uart_tx_inst.n873\ : std_logic;
signal \uart_tx_inst.data_reg_1\ : std_logic;
signal \uart_tx_inst.data_reg_2\ : std_logic;
signal \uart_tx_inst.data_reg_3\ : std_logic;
signal \uart_tx_inst.data_reg_4\ : std_logic;
signal \uart_tx_inst.data_reg_5\ : std_logic;
signal \uart_tx_inst.data_reg_6\ : std_logic;
signal input_axis_tvalid_c : std_logic;
signal \uart_tx_inst.data_reg_8\ : std_logic;
signal \uart_tx_inst.data_reg_7\ : std_logic;
signal \uart_tx_inst.n189\ : std_logic;
signal \uart_tx_inst.data_reg_0\ : std_logic;
signal \uart_tx_inst.n7\ : std_logic;
signal \uart_tx_inst.n15\ : std_logic;
signal txd_c : std_logic;
signal clk_c : std_logic;
signal \uart_tx_inst.n719\ : std_logic;
signal rst_c : std_logic;
signal n108 : std_logic;
signal \bfn_12_5_0_\ : std_logic;
signal n107 : std_logic;
signal \uart_tx_inst.n1582\ : std_logic;
signal n106 : std_logic;
signal \uart_tx_inst.n1583\ : std_logic;
signal n105 : std_logic;
signal \uart_tx_inst.n1584\ : std_logic;
signal n104 : std_logic;
signal \uart_tx_inst.n1585\ : std_logic;
signal n103 : std_logic;
signal \uart_tx_inst.n1586\ : std_logic;
signal n102 : std_logic;
signal \uart_tx_inst.n1587\ : std_logic;
signal n101 : std_logic;
signal \uart_tx_inst.n1588\ : std_logic;
signal \uart_tx_inst.n1589\ : std_logic;
signal input_axis_tdata_c_0 : std_logic;
signal n100 : std_logic;
signal \bfn_12_6_0_\ : std_logic;
signal input_axis_tdata_c_1 : std_logic;
signal n99 : std_logic;
signal \uart_tx_inst.n1590\ : std_logic;
signal input_axis_tdata_c_2 : std_logic;
signal n98 : std_logic;
signal \uart_tx_inst.n1591\ : std_logic;
signal input_axis_tdata_c_3 : std_logic;
signal n97 : std_logic;
signal \uart_tx_inst.n1592\ : std_logic;
signal input_axis_tdata_c_4 : std_logic;
signal n96 : std_logic;
signal \uart_tx_inst.n1593\ : std_logic;
signal input_axis_tdata_c_5 : std_logic;
signal n95 : std_logic;
signal \uart_tx_inst.n1594\ : std_logic;
signal input_axis_tdata_c_6 : std_logic;
signal n94 : std_logic;
signal \uart_tx_inst.n1595\ : std_logic;
signal input_axis_tdata_c_7 : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \uart_tx_inst.n1596\ : std_logic;
signal n93 : std_logic;
signal \_gnd_net_\ : std_logic;

signal clk_wire : std_logic;
signal input_axis_tdata_wire : std_logic_vector(7 downto 0);
signal input_axis_tready_wire : std_logic;
signal input_axis_tvalid_wire : std_logic;
signal output_axis_tdata_wire : std_logic_vector(7 downto 0);
signal output_axis_tready_wire : std_logic;
signal output_axis_tvalid_wire : std_logic;
signal rst_wire : std_logic;
signal rx_busy_wire : std_logic;
signal rx_frame_error_wire : std_logic;
signal rx_overrun_error_wire : std_logic;
signal rxd_wire : std_logic;
signal tx_busy_wire : std_logic;
signal txd_wire : std_logic;

begin
    clk_wire <= clk;
    input_axis_tdata_wire <= input_axis_tdata;
    input_axis_tready <= input_axis_tready_wire;
    input_axis_tvalid_wire <= input_axis_tvalid;
    output_axis_tdata <= output_axis_tdata_wire;
    output_axis_tready_wire <= output_axis_tready;
    output_axis_tvalid <= output_axis_tvalid_wire;
    rst_wire <= rst;
    rx_busy <= rx_busy_wire;
    rx_frame_error <= rx_frame_error_wire;
    rx_overrun_error <= rx_overrun_error_wire;
    rxd_wire <= rxd;
    tx_busy <= tx_busy_wire;
    txd <= txd_wire;

    \clk_pad_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__9134\,
            GLOBALBUFFEROUTPUT => clk_c
        );

    \clk_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9136\,
            DIN => \N__9135\,
            DOUT => \N__9134\,
            PACKAGEPIN => clk_wire
        );

    \clk_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9136\,
            PADOUT => \N__9135\,
            PADIN => \N__9134\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \input_axis_tdata_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9125\,
            DIN => \N__9124\,
            DOUT => \N__9123\,
            PACKAGEPIN => input_axis_tdata_wire(0)
        );

    \input_axis_tdata_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9125\,
            PADOUT => \N__9124\,
            PADIN => \N__9123\,
            CLOCKENABLE => 'H',
            DIN0 => input_axis_tdata_c_0,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \input_axis_tdata_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9116\,
            DIN => \N__9115\,
            DOUT => \N__9114\,
            PACKAGEPIN => input_axis_tdata_wire(1)
        );

    \input_axis_tdata_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9116\,
            PADOUT => \N__9115\,
            PADIN => \N__9114\,
            CLOCKENABLE => 'H',
            DIN0 => input_axis_tdata_c_1,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \input_axis_tdata_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9107\,
            DIN => \N__9106\,
            DOUT => \N__9105\,
            PACKAGEPIN => input_axis_tdata_wire(2)
        );

    \input_axis_tdata_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9107\,
            PADOUT => \N__9106\,
            PADIN => \N__9105\,
            CLOCKENABLE => 'H',
            DIN0 => input_axis_tdata_c_2,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \input_axis_tdata_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9098\,
            DIN => \N__9097\,
            DOUT => \N__9096\,
            PACKAGEPIN => input_axis_tdata_wire(3)
        );

    \input_axis_tdata_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9098\,
            PADOUT => \N__9097\,
            PADIN => \N__9096\,
            CLOCKENABLE => 'H',
            DIN0 => input_axis_tdata_c_3,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \input_axis_tdata_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9089\,
            DIN => \N__9088\,
            DOUT => \N__9087\,
            PACKAGEPIN => input_axis_tdata_wire(4)
        );

    \input_axis_tdata_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9089\,
            PADOUT => \N__9088\,
            PADIN => \N__9087\,
            CLOCKENABLE => 'H',
            DIN0 => input_axis_tdata_c_4,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \input_axis_tdata_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9080\,
            DIN => \N__9079\,
            DOUT => \N__9078\,
            PACKAGEPIN => input_axis_tdata_wire(5)
        );

    \input_axis_tdata_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9080\,
            PADOUT => \N__9079\,
            PADIN => \N__9078\,
            CLOCKENABLE => 'H',
            DIN0 => input_axis_tdata_c_5,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \input_axis_tdata_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9071\,
            DIN => \N__9070\,
            DOUT => \N__9069\,
            PACKAGEPIN => input_axis_tdata_wire(6)
        );

    \input_axis_tdata_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9071\,
            PADOUT => \N__9070\,
            PADIN => \N__9069\,
            CLOCKENABLE => 'H',
            DIN0 => input_axis_tdata_c_6,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \input_axis_tdata_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9062\,
            DIN => \N__9061\,
            DOUT => \N__9060\,
            PACKAGEPIN => input_axis_tdata_wire(7)
        );

    \input_axis_tdata_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9062\,
            PADOUT => \N__9061\,
            PADIN => \N__9060\,
            CLOCKENABLE => 'H',
            DIN0 => input_axis_tdata_c_7,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \input_axis_tready_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9053\,
            DIN => \N__9052\,
            DOUT => \N__9051\,
            PACKAGEPIN => input_axis_tready_wire
        );

    \input_axis_tready_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9053\,
            PADOUT => \N__9052\,
            PADIN => \N__9051\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__3358\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \input_axis_tvalid_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9044\,
            DIN => \N__9043\,
            DOUT => \N__9042\,
            PACKAGEPIN => input_axis_tvalid_wire
        );

    \input_axis_tvalid_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9044\,
            PADOUT => \N__9043\,
            PADIN => \N__9042\,
            CLOCKENABLE => 'H',
            DIN0 => input_axis_tvalid_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \output_axis_tdata_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9035\,
            DIN => \N__9034\,
            DOUT => \N__9033\,
            PACKAGEPIN => output_axis_tdata_wire(0)
        );

    \output_axis_tdata_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9035\,
            PADOUT => \N__9034\,
            PADIN => \N__9033\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__4057\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \output_axis_tdata_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9026\,
            DIN => \N__9025\,
            DOUT => \N__9024\,
            PACKAGEPIN => output_axis_tdata_wire(1)
        );

    \output_axis_tdata_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9026\,
            PADOUT => \N__9025\,
            PADIN => \N__9024\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__5467\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \output_axis_tdata_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9017\,
            DIN => \N__9016\,
            DOUT => \N__9015\,
            PACKAGEPIN => output_axis_tdata_wire(2)
        );

    \output_axis_tdata_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9017\,
            PADOUT => \N__9016\,
            PADIN => \N__9015\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__5137\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \output_axis_tdata_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9008\,
            DIN => \N__9007\,
            DOUT => \N__9006\,
            PACKAGEPIN => output_axis_tdata_wire(3)
        );

    \output_axis_tdata_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9008\,
            PADOUT => \N__9007\,
            PADIN => \N__9006\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__5431\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \output_axis_tdata_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8999\,
            DIN => \N__8998\,
            DOUT => \N__8997\,
            PACKAGEPIN => output_axis_tdata_wire(4)
        );

    \output_axis_tdata_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__8999\,
            PADOUT => \N__8998\,
            PADIN => \N__8997\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__5539\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \output_axis_tdata_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8990\,
            DIN => \N__8989\,
            DOUT => \N__8988\,
            PACKAGEPIN => output_axis_tdata_wire(5)
        );

    \output_axis_tdata_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__8990\,
            PADOUT => \N__8989\,
            PADIN => \N__8988\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__5506\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \output_axis_tdata_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8981\,
            DIN => \N__8980\,
            DOUT => \N__8979\,
            PACKAGEPIN => output_axis_tdata_wire(6)
        );

    \output_axis_tdata_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__8981\,
            PADOUT => \N__8980\,
            PADIN => \N__8979\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__5173\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \output_axis_tdata_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8972\,
            DIN => \N__8971\,
            DOUT => \N__8970\,
            PACKAGEPIN => output_axis_tdata_wire(7)
        );

    \output_axis_tdata_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__8972\,
            PADOUT => \N__8971\,
            PADIN => \N__8970\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__5095\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \output_axis_tready_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8963\,
            DIN => \N__8962\,
            DOUT => \N__8961\,
            PACKAGEPIN => output_axis_tready_wire
        );

    \output_axis_tready_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__8963\,
            PADOUT => \N__8962\,
            PADIN => \N__8961\,
            CLOCKENABLE => 'H',
            DIN0 => output_axis_tready_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \output_axis_tvalid_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8954\,
            DIN => \N__8953\,
            DOUT => \N__8952\,
            PACKAGEPIN => output_axis_tvalid_wire
        );

    \output_axis_tvalid_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__8954\,
            PADOUT => \N__8953\,
            PADIN => \N__8952\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__3607\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rst_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8945\,
            DIN => \N__8944\,
            DOUT => \N__8943\,
            PACKAGEPIN => rst_wire
        );

    \rst_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__8945\,
            PADOUT => \N__8944\,
            PADIN => \N__8943\,
            CLOCKENABLE => 'H',
            DIN0 => rst_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rx_busy_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8936\,
            DIN => \N__8935\,
            DOUT => \N__8934\,
            PACKAGEPIN => rx_busy_wire
        );

    \rx_busy_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__8936\,
            PADOUT => \N__8935\,
            PADIN => \N__8934\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__3322\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rx_frame_error_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8927\,
            DIN => \N__8926\,
            DOUT => \N__8925\,
            PACKAGEPIN => rx_frame_error_wire
        );

    \rx_frame_error_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__8927\,
            PADOUT => \N__8926\,
            PADIN => \N__8925\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__5218\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rx_overrun_error_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8918\,
            DIN => \N__8917\,
            DOUT => \N__8916\,
            PACKAGEPIN => rx_overrun_error_wire
        );

    \rx_overrun_error_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__8918\,
            PADOUT => \N__8917\,
            PADIN => \N__8916\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__3382\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rxd_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8909\,
            DIN => \N__8908\,
            DOUT => \N__8907\,
            PACKAGEPIN => rxd_wire
        );

    \rxd_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__8909\,
            PADOUT => \N__8908\,
            PADIN => \N__8907\,
            CLOCKENABLE => 'H',
            DIN0 => rxd_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \tx_busy_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8900\,
            DIN => \N__8899\,
            DOUT => \N__8898\,
            PACKAGEPIN => tx_busy_wire
        );

    \tx_busy_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__8900\,
            PADOUT => \N__8899\,
            PADIN => \N__8898\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__3304\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \txd_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8891\,
            DIN => \N__8890\,
            DOUT => \N__8889\,
            PACKAGEPIN => txd_wire
        );

    \txd_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__8891\,
            PADOUT => \N__8890\,
            PADIN => \N__8889\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7405\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__2137\ : CascadeMux
    port map (
            O => \N__8872\,
            I => \N__8868\
        );

    \I__2136\ : InMux
    port map (
            O => \N__8871\,
            I => \N__8862\
        );

    \I__2135\ : InMux
    port map (
            O => \N__8868\,
            I => \N__8862\
        );

    \I__2134\ : CascadeMux
    port map (
            O => \N__8867\,
            I => \N__8859\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__8862\,
            I => \N__8855\
        );

    \I__2132\ : InMux
    port map (
            O => \N__8859\,
            I => \N__8852\
        );

    \I__2131\ : CascadeMux
    port map (
            O => \N__8858\,
            I => \N__8849\
        );

    \I__2130\ : Span4Mux_h
    port map (
            O => \N__8855\,
            I => \N__8842\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__8852\,
            I => \N__8842\
        );

    \I__2128\ : InMux
    port map (
            O => \N__8849\,
            I => \N__8839\
        );

    \I__2127\ : CascadeMux
    port map (
            O => \N__8848\,
            I => \N__8836\
        );

    \I__2126\ : CascadeMux
    port map (
            O => \N__8847\,
            I => \N__8832\
        );

    \I__2125\ : Span4Mux_s1_h
    port map (
            O => \N__8842\,
            I => \N__8827\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__8839\,
            I => \N__8827\
        );

    \I__2123\ : InMux
    port map (
            O => \N__8836\,
            I => \N__8824\
        );

    \I__2122\ : CascadeMux
    port map (
            O => \N__8835\,
            I => \N__8821\
        );

    \I__2121\ : InMux
    port map (
            O => \N__8832\,
            I => \N__8818\
        );

    \I__2120\ : Span4Mux_v
    port map (
            O => \N__8827\,
            I => \N__8813\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__8824\,
            I => \N__8813\
        );

    \I__2118\ : InMux
    port map (
            O => \N__8821\,
            I => \N__8810\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__8818\,
            I => input_axis_tdata_c_3
        );

    \I__2116\ : Odrv4
    port map (
            O => \N__8813\,
            I => input_axis_tdata_c_3
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__8810\,
            I => input_axis_tdata_c_3
        );

    \I__2114\ : InMux
    port map (
            O => \N__8803\,
            I => \N__8800\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__8800\,
            I => \N__8796\
        );

    \I__2112\ : InMux
    port map (
            O => \N__8799\,
            I => \N__8793\
        );

    \I__2111\ : Span4Mux_s1_v
    port map (
            O => \N__8796\,
            I => \N__8790\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__8793\,
            I => \N__8787\
        );

    \I__2109\ : Span4Mux_v
    port map (
            O => \N__8790\,
            I => \N__8782\
        );

    \I__2108\ : Span4Mux_v
    port map (
            O => \N__8787\,
            I => \N__8782\
        );

    \I__2107\ : Odrv4
    port map (
            O => \N__8782\,
            I => n97
        );

    \I__2106\ : InMux
    port map (
            O => \N__8779\,
            I => \uart_tx_inst.n1592\
        );

    \I__2105\ : InMux
    port map (
            O => \N__8776\,
            I => \N__8772\
        );

    \I__2104\ : InMux
    port map (
            O => \N__8775\,
            I => \N__8767\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__8772\,
            I => \N__8764\
        );

    \I__2102\ : InMux
    port map (
            O => \N__8771\,
            I => \N__8761\
        );

    \I__2101\ : CascadeMux
    port map (
            O => \N__8770\,
            I => \N__8758\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__8767\,
            I => \N__8754\
        );

    \I__2099\ : Span4Mux_h
    port map (
            O => \N__8764\,
            I => \N__8748\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__8761\,
            I => \N__8748\
        );

    \I__2097\ : InMux
    port map (
            O => \N__8758\,
            I => \N__8745\
        );

    \I__2096\ : CascadeMux
    port map (
            O => \N__8757\,
            I => \N__8742\
        );

    \I__2095\ : Span4Mux_s3_v
    port map (
            O => \N__8754\,
            I => \N__8738\
        );

    \I__2094\ : CascadeMux
    port map (
            O => \N__8753\,
            I => \N__8735\
        );

    \I__2093\ : Span4Mux_s1_h
    port map (
            O => \N__8748\,
            I => \N__8730\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__8745\,
            I => \N__8730\
        );

    \I__2091\ : InMux
    port map (
            O => \N__8742\,
            I => \N__8727\
        );

    \I__2090\ : CascadeMux
    port map (
            O => \N__8741\,
            I => \N__8724\
        );

    \I__2089\ : IoSpan4Mux
    port map (
            O => \N__8738\,
            I => \N__8721\
        );

    \I__2088\ : InMux
    port map (
            O => \N__8735\,
            I => \N__8718\
        );

    \I__2087\ : Span4Mux_v
    port map (
            O => \N__8730\,
            I => \N__8713\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__8727\,
            I => \N__8713\
        );

    \I__2085\ : InMux
    port map (
            O => \N__8724\,
            I => \N__8710\
        );

    \I__2084\ : Odrv4
    port map (
            O => \N__8721\,
            I => input_axis_tdata_c_4
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__8718\,
            I => input_axis_tdata_c_4
        );

    \I__2082\ : Odrv4
    port map (
            O => \N__8713\,
            I => input_axis_tdata_c_4
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__8710\,
            I => input_axis_tdata_c_4
        );

    \I__2080\ : InMux
    port map (
            O => \N__8701\,
            I => \N__8698\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__8698\,
            I => \N__8694\
        );

    \I__2078\ : InMux
    port map (
            O => \N__8697\,
            I => \N__8691\
        );

    \I__2077\ : Span4Mux_s1_v
    port map (
            O => \N__8694\,
            I => \N__8688\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__8691\,
            I => \N__8685\
        );

    \I__2075\ : Span4Mux_v
    port map (
            O => \N__8688\,
            I => \N__8680\
        );

    \I__2074\ : Span4Mux_v
    port map (
            O => \N__8685\,
            I => \N__8680\
        );

    \I__2073\ : Odrv4
    port map (
            O => \N__8680\,
            I => n96
        );

    \I__2072\ : InMux
    port map (
            O => \N__8677\,
            I => \uart_tx_inst.n1593\
        );

    \I__2071\ : CascadeMux
    port map (
            O => \N__8674\,
            I => \N__8670\
        );

    \I__2070\ : CascadeMux
    port map (
            O => \N__8673\,
            I => \N__8664\
        );

    \I__2069\ : InMux
    port map (
            O => \N__8670\,
            I => \N__8660\
        );

    \I__2068\ : CascadeMux
    port map (
            O => \N__8669\,
            I => \N__8657\
        );

    \I__2067\ : CascadeMux
    port map (
            O => \N__8668\,
            I => \N__8654\
        );

    \I__2066\ : InMux
    port map (
            O => \N__8667\,
            I => \N__8651\
        );

    \I__2065\ : InMux
    port map (
            O => \N__8664\,
            I => \N__8648\
        );

    \I__2064\ : CascadeMux
    port map (
            O => \N__8663\,
            I => \N__8645\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__8660\,
            I => \N__8642\
        );

    \I__2062\ : InMux
    port map (
            O => \N__8657\,
            I => \N__8639\
        );

    \I__2061\ : InMux
    port map (
            O => \N__8654\,
            I => \N__8636\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__8651\,
            I => \N__8633\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__8648\,
            I => \N__8630\
        );

    \I__2058\ : InMux
    port map (
            O => \N__8645\,
            I => \N__8627\
        );

    \I__2057\ : Span4Mux_h
    port map (
            O => \N__8642\,
            I => \N__8619\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__8639\,
            I => \N__8619\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__8636\,
            I => \N__8619\
        );

    \I__2054\ : Span4Mux_s2_v
    port map (
            O => \N__8633\,
            I => \N__8612\
        );

    \I__2053\ : Span4Mux_s2_v
    port map (
            O => \N__8630\,
            I => \N__8612\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__8627\,
            I => \N__8612\
        );

    \I__2051\ : CascadeMux
    port map (
            O => \N__8626\,
            I => \N__8609\
        );

    \I__2050\ : Span4Mux_v
    port map (
            O => \N__8619\,
            I => \N__8604\
        );

    \I__2049\ : Span4Mux_v
    port map (
            O => \N__8612\,
            I => \N__8604\
        );

    \I__2048\ : InMux
    port map (
            O => \N__8609\,
            I => \N__8601\
        );

    \I__2047\ : Odrv4
    port map (
            O => \N__8604\,
            I => input_axis_tdata_c_5
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__8601\,
            I => input_axis_tdata_c_5
        );

    \I__2045\ : InMux
    port map (
            O => \N__8596\,
            I => \N__8592\
        );

    \I__2044\ : InMux
    port map (
            O => \N__8595\,
            I => \N__8589\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__8592\,
            I => \N__8586\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__8589\,
            I => \N__8583\
        );

    \I__2041\ : Span4Mux_v
    port map (
            O => \N__8586\,
            I => \N__8578\
        );

    \I__2040\ : Span4Mux_v
    port map (
            O => \N__8583\,
            I => \N__8578\
        );

    \I__2039\ : Odrv4
    port map (
            O => \N__8578\,
            I => n95
        );

    \I__2038\ : InMux
    port map (
            O => \N__8575\,
            I => \uart_tx_inst.n1594\
        );

    \I__2037\ : CascadeMux
    port map (
            O => \N__8572\,
            I => \N__8567\
        );

    \I__2036\ : InMux
    port map (
            O => \N__8571\,
            I => \N__8561\
        );

    \I__2035\ : InMux
    port map (
            O => \N__8570\,
            I => \N__8558\
        );

    \I__2034\ : InMux
    port map (
            O => \N__8567\,
            I => \N__8555\
        );

    \I__2033\ : CascadeMux
    port map (
            O => \N__8566\,
            I => \N__8552\
        );

    \I__2032\ : CascadeMux
    port map (
            O => \N__8565\,
            I => \N__8549\
        );

    \I__2031\ : CascadeMux
    port map (
            O => \N__8564\,
            I => \N__8546\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__8561\,
            I => \N__8543\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__8558\,
            I => \N__8538\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__8555\,
            I => \N__8538\
        );

    \I__2027\ : InMux
    port map (
            O => \N__8552\,
            I => \N__8535\
        );

    \I__2026\ : InMux
    port map (
            O => \N__8549\,
            I => \N__8532\
        );

    \I__2025\ : InMux
    port map (
            O => \N__8546\,
            I => \N__8529\
        );

    \I__2024\ : Span4Mux_s2_v
    port map (
            O => \N__8543\,
            I => \N__8525\
        );

    \I__2023\ : Span4Mux_s2_v
    port map (
            O => \N__8538\,
            I => \N__8518\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__8535\,
            I => \N__8518\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__8532\,
            I => \N__8518\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__8529\,
            I => \N__8515\
        );

    \I__2019\ : CascadeMux
    port map (
            O => \N__8528\,
            I => \N__8512\
        );

    \I__2018\ : Span4Mux_v
    port map (
            O => \N__8525\,
            I => \N__8509\
        );

    \I__2017\ : Span4Mux_v
    port map (
            O => \N__8518\,
            I => \N__8506\
        );

    \I__2016\ : Span4Mux_v
    port map (
            O => \N__8515\,
            I => \N__8503\
        );

    \I__2015\ : InMux
    port map (
            O => \N__8512\,
            I => \N__8500\
        );

    \I__2014\ : Odrv4
    port map (
            O => \N__8509\,
            I => input_axis_tdata_c_6
        );

    \I__2013\ : Odrv4
    port map (
            O => \N__8506\,
            I => input_axis_tdata_c_6
        );

    \I__2012\ : Odrv4
    port map (
            O => \N__8503\,
            I => input_axis_tdata_c_6
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__8500\,
            I => input_axis_tdata_c_6
        );

    \I__2010\ : InMux
    port map (
            O => \N__8491\,
            I => \N__8488\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__8488\,
            I => \N__8484\
        );

    \I__2008\ : InMux
    port map (
            O => \N__8487\,
            I => \N__8481\
        );

    \I__2007\ : Span4Mux_s1_v
    port map (
            O => \N__8484\,
            I => \N__8478\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__8481\,
            I => \N__8475\
        );

    \I__2005\ : Span4Mux_v
    port map (
            O => \N__8478\,
            I => \N__8470\
        );

    \I__2004\ : Span4Mux_v
    port map (
            O => \N__8475\,
            I => \N__8470\
        );

    \I__2003\ : Odrv4
    port map (
            O => \N__8470\,
            I => n94
        );

    \I__2002\ : InMux
    port map (
            O => \N__8467\,
            I => \uart_tx_inst.n1595\
        );

    \I__2001\ : CascadeMux
    port map (
            O => \N__8464\,
            I => \N__8459\
        );

    \I__2000\ : CascadeMux
    port map (
            O => \N__8463\,
            I => \N__8455\
        );

    \I__1999\ : InMux
    port map (
            O => \N__8462\,
            I => \N__8450\
        );

    \I__1998\ : InMux
    port map (
            O => \N__8459\,
            I => \N__8447\
        );

    \I__1997\ : CascadeMux
    port map (
            O => \N__8458\,
            I => \N__8444\
        );

    \I__1996\ : InMux
    port map (
            O => \N__8455\,
            I => \N__8441\
        );

    \I__1995\ : CascadeMux
    port map (
            O => \N__8454\,
            I => \N__8438\
        );

    \I__1994\ : CascadeMux
    port map (
            O => \N__8453\,
            I => \N__8435\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__8450\,
            I => \N__8429\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__8447\,
            I => \N__8429\
        );

    \I__1991\ : InMux
    port map (
            O => \N__8444\,
            I => \N__8426\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__8441\,
            I => \N__8423\
        );

    \I__1989\ : InMux
    port map (
            O => \N__8438\,
            I => \N__8420\
        );

    \I__1988\ : InMux
    port map (
            O => \N__8435\,
            I => \N__8417\
        );

    \I__1987\ : InMux
    port map (
            O => \N__8434\,
            I => \N__8414\
        );

    \I__1986\ : Span4Mux_s3_v
    port map (
            O => \N__8429\,
            I => \N__8411\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__8426\,
            I => \N__8404\
        );

    \I__1984\ : Sp12to4
    port map (
            O => \N__8423\,
            I => \N__8404\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__8420\,
            I => \N__8404\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__8417\,
            I => \N__8399\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__8414\,
            I => \N__8399\
        );

    \I__1980\ : Span4Mux_v
    port map (
            O => \N__8411\,
            I => \N__8396\
        );

    \I__1979\ : Span12Mux_s7_v
    port map (
            O => \N__8404\,
            I => \N__8393\
        );

    \I__1978\ : Span4Mux_v
    port map (
            O => \N__8399\,
            I => \N__8390\
        );

    \I__1977\ : Odrv4
    port map (
            O => \N__8396\,
            I => input_axis_tdata_c_7
        );

    \I__1976\ : Odrv12
    port map (
            O => \N__8393\,
            I => input_axis_tdata_c_7
        );

    \I__1975\ : Odrv4
    port map (
            O => \N__8390\,
            I => input_axis_tdata_c_7
        );

    \I__1974\ : CascadeMux
    port map (
            O => \N__8383\,
            I => \N__8371\
        );

    \I__1973\ : CascadeMux
    port map (
            O => \N__8382\,
            I => \N__8367\
        );

    \I__1972\ : CascadeMux
    port map (
            O => \N__8381\,
            I => \N__8363\
        );

    \I__1971\ : CascadeMux
    port map (
            O => \N__8380\,
            I => \N__8360\
        );

    \I__1970\ : CascadeMux
    port map (
            O => \N__8379\,
            I => \N__8356\
        );

    \I__1969\ : CascadeMux
    port map (
            O => \N__8378\,
            I => \N__8352\
        );

    \I__1968\ : CascadeMux
    port map (
            O => \N__8377\,
            I => \N__8348\
        );

    \I__1967\ : CascadeMux
    port map (
            O => \N__8376\,
            I => \N__8344\
        );

    \I__1966\ : CascadeMux
    port map (
            O => \N__8375\,
            I => \N__8339\
        );

    \I__1965\ : CascadeMux
    port map (
            O => \N__8374\,
            I => \N__8336\
        );

    \I__1964\ : InMux
    port map (
            O => \N__8371\,
            I => \N__8315\
        );

    \I__1963\ : InMux
    port map (
            O => \N__8370\,
            I => \N__8315\
        );

    \I__1962\ : InMux
    port map (
            O => \N__8367\,
            I => \N__8315\
        );

    \I__1961\ : InMux
    port map (
            O => \N__8366\,
            I => \N__8315\
        );

    \I__1960\ : InMux
    port map (
            O => \N__8363\,
            I => \N__8315\
        );

    \I__1959\ : InMux
    port map (
            O => \N__8360\,
            I => \N__8315\
        );

    \I__1958\ : InMux
    port map (
            O => \N__8359\,
            I => \N__8298\
        );

    \I__1957\ : InMux
    port map (
            O => \N__8356\,
            I => \N__8298\
        );

    \I__1956\ : InMux
    port map (
            O => \N__8355\,
            I => \N__8298\
        );

    \I__1955\ : InMux
    port map (
            O => \N__8352\,
            I => \N__8298\
        );

    \I__1954\ : InMux
    port map (
            O => \N__8351\,
            I => \N__8298\
        );

    \I__1953\ : InMux
    port map (
            O => \N__8348\,
            I => \N__8298\
        );

    \I__1952\ : InMux
    port map (
            O => \N__8347\,
            I => \N__8298\
        );

    \I__1951\ : InMux
    port map (
            O => \N__8344\,
            I => \N__8298\
        );

    \I__1950\ : InMux
    port map (
            O => \N__8343\,
            I => \N__8291\
        );

    \I__1949\ : InMux
    port map (
            O => \N__8342\,
            I => \N__8291\
        );

    \I__1948\ : InMux
    port map (
            O => \N__8339\,
            I => \N__8291\
        );

    \I__1947\ : InMux
    port map (
            O => \N__8336\,
            I => \N__8288\
        );

    \I__1946\ : InMux
    port map (
            O => \N__8335\,
            I => \N__8279\
        );

    \I__1945\ : InMux
    port map (
            O => \N__8334\,
            I => \N__8279\
        );

    \I__1944\ : InMux
    port map (
            O => \N__8333\,
            I => \N__8279\
        );

    \I__1943\ : InMux
    port map (
            O => \N__8332\,
            I => \N__8279\
        );

    \I__1942\ : InMux
    port map (
            O => \N__8331\,
            I => \N__8270\
        );

    \I__1941\ : InMux
    port map (
            O => \N__8330\,
            I => \N__8270\
        );

    \I__1940\ : InMux
    port map (
            O => \N__8329\,
            I => \N__8270\
        );

    \I__1939\ : InMux
    port map (
            O => \N__8328\,
            I => \N__8270\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__8315\,
            I => \N__8248\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__8298\,
            I => \N__8248\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__8291\,
            I => \N__8248\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__8288\,
            I => \N__8238\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__8279\,
            I => \N__8233\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__8270\,
            I => \N__8233\
        );

    \I__1932\ : InMux
    port map (
            O => \N__8269\,
            I => \N__8224\
        );

    \I__1931\ : InMux
    port map (
            O => \N__8268\,
            I => \N__8224\
        );

    \I__1930\ : InMux
    port map (
            O => \N__8267\,
            I => \N__8224\
        );

    \I__1929\ : InMux
    port map (
            O => \N__8266\,
            I => \N__8224\
        );

    \I__1928\ : InMux
    port map (
            O => \N__8265\,
            I => \N__8215\
        );

    \I__1927\ : InMux
    port map (
            O => \N__8264\,
            I => \N__8215\
        );

    \I__1926\ : InMux
    port map (
            O => \N__8263\,
            I => \N__8215\
        );

    \I__1925\ : InMux
    port map (
            O => \N__8262\,
            I => \N__8215\
        );

    \I__1924\ : InMux
    port map (
            O => \N__8261\,
            I => \N__8208\
        );

    \I__1923\ : InMux
    port map (
            O => \N__8260\,
            I => \N__8208\
        );

    \I__1922\ : InMux
    port map (
            O => \N__8259\,
            I => \N__8208\
        );

    \I__1921\ : InMux
    port map (
            O => \N__8258\,
            I => \N__8199\
        );

    \I__1920\ : InMux
    port map (
            O => \N__8257\,
            I => \N__8199\
        );

    \I__1919\ : InMux
    port map (
            O => \N__8256\,
            I => \N__8199\
        );

    \I__1918\ : InMux
    port map (
            O => \N__8255\,
            I => \N__8199\
        );

    \I__1917\ : Span4Mux_v
    port map (
            O => \N__8248\,
            I => \N__8196\
        );

    \I__1916\ : InMux
    port map (
            O => \N__8247\,
            I => \N__8189\
        );

    \I__1915\ : InMux
    port map (
            O => \N__8246\,
            I => \N__8189\
        );

    \I__1914\ : InMux
    port map (
            O => \N__8245\,
            I => \N__8189\
        );

    \I__1913\ : InMux
    port map (
            O => \N__8244\,
            I => \N__8180\
        );

    \I__1912\ : InMux
    port map (
            O => \N__8243\,
            I => \N__8180\
        );

    \I__1911\ : InMux
    port map (
            O => \N__8242\,
            I => \N__8180\
        );

    \I__1910\ : InMux
    port map (
            O => \N__8241\,
            I => \N__8180\
        );

    \I__1909\ : Span4Mux_s2_h
    port map (
            O => \N__8238\,
            I => \N__8175\
        );

    \I__1908\ : Span4Mux_s2_h
    port map (
            O => \N__8233\,
            I => \N__8175\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__8224\,
            I => \N__8170\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__8215\,
            I => \N__8170\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__8208\,
            I => \N__8158\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__8199\,
            I => \N__8158\
        );

    \I__1903\ : Sp12to4
    port map (
            O => \N__8196\,
            I => \N__8158\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__8189\,
            I => \N__8158\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__8180\,
            I => \N__8158\
        );

    \I__1900\ : Span4Mux_v
    port map (
            O => \N__8175\,
            I => \N__8153\
        );

    \I__1899\ : Span4Mux_s2_h
    port map (
            O => \N__8170\,
            I => \N__8153\
        );

    \I__1898\ : InMux
    port map (
            O => \N__8169\,
            I => \N__8150\
        );

    \I__1897\ : Span12Mux_s6_h
    port map (
            O => \N__8158\,
            I => \N__8147\
        );

    \I__1896\ : Span4Mux_h
    port map (
            O => \N__8153\,
            I => \N__8144\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__8150\,
            I => \N__8141\
        );

    \I__1894\ : Odrv12
    port map (
            O => \N__8147\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1893\ : Odrv4
    port map (
            O => \N__8144\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1892\ : Odrv12
    port map (
            O => \N__8141\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1891\ : InMux
    port map (
            O => \N__8134\,
            I => \uart_tx_inst.n1596\
        );

    \I__1890\ : InMux
    port map (
            O => \N__8131\,
            I => \N__8127\
        );

    \I__1889\ : InMux
    port map (
            O => \N__8130\,
            I => \N__8124\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__8127\,
            I => \N__8121\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__8124\,
            I => \N__8118\
        );

    \I__1886\ : Span4Mux_v
    port map (
            O => \N__8121\,
            I => \N__8113\
        );

    \I__1885\ : Span4Mux_v
    port map (
            O => \N__8118\,
            I => \N__8113\
        );

    \I__1884\ : Odrv4
    port map (
            O => \N__8113\,
            I => n93
        );

    \I__1883\ : InMux
    port map (
            O => \N__8110\,
            I => \uart_tx_inst.n1583\
        );

    \I__1882\ : InMux
    port map (
            O => \N__8107\,
            I => \N__8103\
        );

    \I__1881\ : InMux
    port map (
            O => \N__8106\,
            I => \N__8100\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__8103\,
            I => \N__8097\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__8100\,
            I => \N__8094\
        );

    \I__1878\ : Span4Mux_h
    port map (
            O => \N__8097\,
            I => \N__8091\
        );

    \I__1877\ : Span4Mux_h
    port map (
            O => \N__8094\,
            I => \N__8088\
        );

    \I__1876\ : Odrv4
    port map (
            O => \N__8091\,
            I => n105
        );

    \I__1875\ : Odrv4
    port map (
            O => \N__8088\,
            I => n105
        );

    \I__1874\ : InMux
    port map (
            O => \N__8083\,
            I => \uart_tx_inst.n1584\
        );

    \I__1873\ : InMux
    port map (
            O => \N__8080\,
            I => \N__8076\
        );

    \I__1872\ : InMux
    port map (
            O => \N__8079\,
            I => \N__8073\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__8076\,
            I => \N__8070\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__8073\,
            I => \N__8067\
        );

    \I__1869\ : Span4Mux_v
    port map (
            O => \N__8070\,
            I => \N__8062\
        );

    \I__1868\ : Span4Mux_v
    port map (
            O => \N__8067\,
            I => \N__8062\
        );

    \I__1867\ : Odrv4
    port map (
            O => \N__8062\,
            I => n104
        );

    \I__1866\ : InMux
    port map (
            O => \N__8059\,
            I => \uart_tx_inst.n1585\
        );

    \I__1865\ : InMux
    port map (
            O => \N__8056\,
            I => \N__8052\
        );

    \I__1864\ : InMux
    port map (
            O => \N__8055\,
            I => \N__8049\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__8052\,
            I => \N__8046\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__8049\,
            I => \N__8043\
        );

    \I__1861\ : Span4Mux_v
    port map (
            O => \N__8046\,
            I => \N__8040\
        );

    \I__1860\ : Span4Mux_s3_v
    port map (
            O => \N__8043\,
            I => \N__8037\
        );

    \I__1859\ : Odrv4
    port map (
            O => \N__8040\,
            I => n103
        );

    \I__1858\ : Odrv4
    port map (
            O => \N__8037\,
            I => n103
        );

    \I__1857\ : InMux
    port map (
            O => \N__8032\,
            I => \uart_tx_inst.n1586\
        );

    \I__1856\ : InMux
    port map (
            O => \N__8029\,
            I => \N__8025\
        );

    \I__1855\ : InMux
    port map (
            O => \N__8028\,
            I => \N__8022\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__8025\,
            I => \N__8019\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__8022\,
            I => \N__8016\
        );

    \I__1852\ : Span4Mux_s3_v
    port map (
            O => \N__8019\,
            I => \N__8013\
        );

    \I__1851\ : Span4Mux_v
    port map (
            O => \N__8016\,
            I => \N__8010\
        );

    \I__1850\ : Odrv4
    port map (
            O => \N__8013\,
            I => n102
        );

    \I__1849\ : Odrv4
    port map (
            O => \N__8010\,
            I => n102
        );

    \I__1848\ : InMux
    port map (
            O => \N__8005\,
            I => \uart_tx_inst.n1587\
        );

    \I__1847\ : InMux
    port map (
            O => \N__8002\,
            I => \N__7999\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__7999\,
            I => \N__7995\
        );

    \I__1845\ : InMux
    port map (
            O => \N__7998\,
            I => \N__7992\
        );

    \I__1844\ : Span4Mux_v
    port map (
            O => \N__7995\,
            I => \N__7989\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__7992\,
            I => \N__7986\
        );

    \I__1842\ : Span4Mux_h
    port map (
            O => \N__7989\,
            I => \N__7983\
        );

    \I__1841\ : Span12Mux_s4_v
    port map (
            O => \N__7986\,
            I => \N__7980\
        );

    \I__1840\ : Odrv4
    port map (
            O => \N__7983\,
            I => n101
        );

    \I__1839\ : Odrv12
    port map (
            O => \N__7980\,
            I => n101
        );

    \I__1838\ : InMux
    port map (
            O => \N__7975\,
            I => \uart_tx_inst.n1588\
        );

    \I__1837\ : CascadeMux
    port map (
            O => \N__7972\,
            I => \N__7966\
        );

    \I__1836\ : CascadeMux
    port map (
            O => \N__7971\,
            I => \N__7963\
        );

    \I__1835\ : InMux
    port map (
            O => \N__7970\,
            I => \N__7960\
        );

    \I__1834\ : InMux
    port map (
            O => \N__7969\,
            I => \N__7955\
        );

    \I__1833\ : InMux
    port map (
            O => \N__7966\,
            I => \N__7952\
        );

    \I__1832\ : InMux
    port map (
            O => \N__7963\,
            I => \N__7949\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__7960\,
            I => \N__7946\
        );

    \I__1830\ : InMux
    port map (
            O => \N__7959\,
            I => \N__7943\
        );

    \I__1829\ : InMux
    port map (
            O => \N__7958\,
            I => \N__7940\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__7955\,
            I => \N__7936\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__7952\,
            I => \N__7925\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__7949\,
            I => \N__7925\
        );

    \I__1825\ : Span4Mux_s2_v
    port map (
            O => \N__7946\,
            I => \N__7925\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__7943\,
            I => \N__7925\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__7940\,
            I => \N__7925\
        );

    \I__1822\ : CascadeMux
    port map (
            O => \N__7939\,
            I => \N__7922\
        );

    \I__1821\ : Span4Mux_h
    port map (
            O => \N__7936\,
            I => \N__7917\
        );

    \I__1820\ : Span4Mux_v
    port map (
            O => \N__7925\,
            I => \N__7917\
        );

    \I__1819\ : InMux
    port map (
            O => \N__7922\,
            I => \N__7914\
        );

    \I__1818\ : Odrv4
    port map (
            O => \N__7917\,
            I => input_axis_tdata_c_0
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__7914\,
            I => input_axis_tdata_c_0
        );

    \I__1816\ : InMux
    port map (
            O => \N__7909\,
            I => \N__7906\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__7906\,
            I => \N__7902\
        );

    \I__1814\ : InMux
    port map (
            O => \N__7905\,
            I => \N__7899\
        );

    \I__1813\ : Span4Mux_v
    port map (
            O => \N__7902\,
            I => \N__7894\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__7899\,
            I => \N__7894\
        );

    \I__1811\ : Span4Mux_v
    port map (
            O => \N__7894\,
            I => \N__7891\
        );

    \I__1810\ : Odrv4
    port map (
            O => \N__7891\,
            I => n100
        );

    \I__1809\ : InMux
    port map (
            O => \N__7888\,
            I => \bfn_12_6_0_\
        );

    \I__1808\ : CascadeMux
    port map (
            O => \N__7885\,
            I => \N__7878\
        );

    \I__1807\ : CascadeMux
    port map (
            O => \N__7884\,
            I => \N__7874\
        );

    \I__1806\ : InMux
    port map (
            O => \N__7883\,
            I => \N__7871\
        );

    \I__1805\ : CascadeMux
    port map (
            O => \N__7882\,
            I => \N__7868\
        );

    \I__1804\ : CascadeMux
    port map (
            O => \N__7881\,
            I => \N__7865\
        );

    \I__1803\ : InMux
    port map (
            O => \N__7878\,
            I => \N__7862\
        );

    \I__1802\ : InMux
    port map (
            O => \N__7877\,
            I => \N__7859\
        );

    \I__1801\ : InMux
    port map (
            O => \N__7874\,
            I => \N__7856\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__7871\,
            I => \N__7853\
        );

    \I__1799\ : InMux
    port map (
            O => \N__7868\,
            I => \N__7850\
        );

    \I__1798\ : InMux
    port map (
            O => \N__7865\,
            I => \N__7847\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__7862\,
            I => \N__7843\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__7859\,
            I => \N__7838\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__7856\,
            I => \N__7838\
        );

    \I__1794\ : Span4Mux_s3_v
    port map (
            O => \N__7853\,
            I => \N__7831\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__7850\,
            I => \N__7831\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__7847\,
            I => \N__7831\
        );

    \I__1791\ : CascadeMux
    port map (
            O => \N__7846\,
            I => \N__7828\
        );

    \I__1790\ : Span4Mux_v
    port map (
            O => \N__7843\,
            I => \N__7821\
        );

    \I__1789\ : Span4Mux_s3_v
    port map (
            O => \N__7838\,
            I => \N__7821\
        );

    \I__1788\ : Span4Mux_v
    port map (
            O => \N__7831\,
            I => \N__7821\
        );

    \I__1787\ : InMux
    port map (
            O => \N__7828\,
            I => \N__7818\
        );

    \I__1786\ : Odrv4
    port map (
            O => \N__7821\,
            I => input_axis_tdata_c_1
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__7818\,
            I => input_axis_tdata_c_1
        );

    \I__1784\ : InMux
    port map (
            O => \N__7813\,
            I => \N__7810\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__7810\,
            I => \N__7806\
        );

    \I__1782\ : InMux
    port map (
            O => \N__7809\,
            I => \N__7803\
        );

    \I__1781\ : Span4Mux_s2_v
    port map (
            O => \N__7806\,
            I => \N__7800\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__7803\,
            I => \N__7797\
        );

    \I__1779\ : Odrv4
    port map (
            O => \N__7800\,
            I => n99
        );

    \I__1778\ : Odrv4
    port map (
            O => \N__7797\,
            I => n99
        );

    \I__1777\ : InMux
    port map (
            O => \N__7792\,
            I => \uart_tx_inst.n1590\
        );

    \I__1776\ : CascadeMux
    port map (
            O => \N__7789\,
            I => \N__7781\
        );

    \I__1775\ : InMux
    port map (
            O => \N__7788\,
            I => \N__7778\
        );

    \I__1774\ : CascadeMux
    port map (
            O => \N__7787\,
            I => \N__7775\
        );

    \I__1773\ : CascadeMux
    port map (
            O => \N__7786\,
            I => \N__7772\
        );

    \I__1772\ : CascadeMux
    port map (
            O => \N__7785\,
            I => \N__7769\
        );

    \I__1771\ : InMux
    port map (
            O => \N__7784\,
            I => \N__7766\
        );

    \I__1770\ : InMux
    port map (
            O => \N__7781\,
            I => \N__7763\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__7778\,
            I => \N__7760\
        );

    \I__1768\ : InMux
    port map (
            O => \N__7775\,
            I => \N__7757\
        );

    \I__1767\ : InMux
    port map (
            O => \N__7772\,
            I => \N__7754\
        );

    \I__1766\ : InMux
    port map (
            O => \N__7769\,
            I => \N__7751\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__7766\,
            I => \N__7747\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__7763\,
            I => \N__7744\
        );

    \I__1763\ : Span4Mux_s3_v
    port map (
            O => \N__7760\,
            I => \N__7735\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__7757\,
            I => \N__7735\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__7754\,
            I => \N__7735\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__7751\,
            I => \N__7735\
        );

    \I__1759\ : CascadeMux
    port map (
            O => \N__7750\,
            I => \N__7732\
        );

    \I__1758\ : IoSpan4Mux
    port map (
            O => \N__7747\,
            I => \N__7729\
        );

    \I__1757\ : Span4Mux_s3_v
    port map (
            O => \N__7744\,
            I => \N__7724\
        );

    \I__1756\ : Span4Mux_v
    port map (
            O => \N__7735\,
            I => \N__7724\
        );

    \I__1755\ : InMux
    port map (
            O => \N__7732\,
            I => \N__7721\
        );

    \I__1754\ : Odrv4
    port map (
            O => \N__7729\,
            I => input_axis_tdata_c_2
        );

    \I__1753\ : Odrv4
    port map (
            O => \N__7724\,
            I => input_axis_tdata_c_2
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__7721\,
            I => input_axis_tdata_c_2
        );

    \I__1751\ : InMux
    port map (
            O => \N__7714\,
            I => \N__7711\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__7711\,
            I => \N__7708\
        );

    \I__1749\ : Span4Mux_s1_v
    port map (
            O => \N__7708\,
            I => \N__7704\
        );

    \I__1748\ : InMux
    port map (
            O => \N__7707\,
            I => \N__7701\
        );

    \I__1747\ : Span4Mux_v
    port map (
            O => \N__7704\,
            I => \N__7696\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__7701\,
            I => \N__7696\
        );

    \I__1745\ : Span4Mux_v
    port map (
            O => \N__7696\,
            I => \N__7693\
        );

    \I__1744\ : Odrv4
    port map (
            O => \N__7693\,
            I => n98
        );

    \I__1743\ : InMux
    port map (
            O => \N__7690\,
            I => \uart_tx_inst.n1591\
        );

    \I__1742\ : InMux
    port map (
            O => \N__7687\,
            I => \N__7684\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__7684\,
            I => \uart_tx_inst.data_reg_3\
        );

    \I__1740\ : InMux
    port map (
            O => \N__7681\,
            I => \N__7678\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__7678\,
            I => \uart_tx_inst.data_reg_4\
        );

    \I__1738\ : CascadeMux
    port map (
            O => \N__7675\,
            I => \N__7672\
        );

    \I__1737\ : InMux
    port map (
            O => \N__7672\,
            I => \N__7669\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__7669\,
            I => \uart_tx_inst.data_reg_5\
        );

    \I__1735\ : InMux
    port map (
            O => \N__7666\,
            I => \N__7663\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__7663\,
            I => \uart_tx_inst.data_reg_6\
        );

    \I__1733\ : InMux
    port map (
            O => \N__7660\,
            I => \N__7646\
        );

    \I__1732\ : CascadeMux
    port map (
            O => \N__7659\,
            I => \N__7642\
        );

    \I__1731\ : CascadeMux
    port map (
            O => \N__7658\,
            I => \N__7639\
        );

    \I__1730\ : InMux
    port map (
            O => \N__7657\,
            I => \N__7622\
        );

    \I__1729\ : InMux
    port map (
            O => \N__7656\,
            I => \N__7622\
        );

    \I__1728\ : InMux
    port map (
            O => \N__7655\,
            I => \N__7622\
        );

    \I__1727\ : InMux
    port map (
            O => \N__7654\,
            I => \N__7622\
        );

    \I__1726\ : InMux
    port map (
            O => \N__7653\,
            I => \N__7622\
        );

    \I__1725\ : InMux
    port map (
            O => \N__7652\,
            I => \N__7622\
        );

    \I__1724\ : InMux
    port map (
            O => \N__7651\,
            I => \N__7622\
        );

    \I__1723\ : InMux
    port map (
            O => \N__7650\,
            I => \N__7622\
        );

    \I__1722\ : InMux
    port map (
            O => \N__7649\,
            I => \N__7619\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__7646\,
            I => \N__7616\
        );

    \I__1720\ : InMux
    port map (
            O => \N__7645\,
            I => \N__7613\
        );

    \I__1719\ : InMux
    port map (
            O => \N__7642\,
            I => \N__7608\
        );

    \I__1718\ : InMux
    port map (
            O => \N__7639\,
            I => \N__7608\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__7622\,
            I => \N__7602\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__7619\,
            I => \N__7595\
        );

    \I__1715\ : Span4Mux_s1_v
    port map (
            O => \N__7616\,
            I => \N__7595\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__7613\,
            I => \N__7595\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__7608\,
            I => \N__7592\
        );

    \I__1712\ : InMux
    port map (
            O => \N__7607\,
            I => \N__7585\
        );

    \I__1711\ : InMux
    port map (
            O => \N__7606\,
            I => \N__7585\
        );

    \I__1710\ : InMux
    port map (
            O => \N__7605\,
            I => \N__7585\
        );

    \I__1709\ : Span4Mux_s3_h
    port map (
            O => \N__7602\,
            I => \N__7580\
        );

    \I__1708\ : Span4Mux_h
    port map (
            O => \N__7595\,
            I => \N__7580\
        );

    \I__1707\ : Span4Mux_h
    port map (
            O => \N__7592\,
            I => \N__7575\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__7585\,
            I => \N__7575\
        );

    \I__1705\ : Odrv4
    port map (
            O => \N__7580\,
            I => input_axis_tvalid_c
        );

    \I__1704\ : Odrv4
    port map (
            O => \N__7575\,
            I => input_axis_tvalid_c
        );

    \I__1703\ : InMux
    port map (
            O => \N__7570\,
            I => \N__7567\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__7567\,
            I => \N__7564\
        );

    \I__1701\ : Span4Mux_s0_h
    port map (
            O => \N__7564\,
            I => \N__7560\
        );

    \I__1700\ : InMux
    port map (
            O => \N__7563\,
            I => \N__7557\
        );

    \I__1699\ : Odrv4
    port map (
            O => \N__7560\,
            I => \uart_tx_inst.data_reg_8\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__7557\,
            I => \uart_tx_inst.data_reg_8\
        );

    \I__1697\ : InMux
    port map (
            O => \N__7552\,
            I => \N__7549\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__7549\,
            I => \uart_tx_inst.data_reg_7\
        );

    \I__1695\ : CEMux
    port map (
            O => \N__7546\,
            I => \N__7543\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__7543\,
            I => \N__7540\
        );

    \I__1693\ : Span4Mux_s0_h
    port map (
            O => \N__7540\,
            I => \N__7537\
        );

    \I__1692\ : Odrv4
    port map (
            O => \N__7537\,
            I => \uart_tx_inst.n189\
        );

    \I__1691\ : InMux
    port map (
            O => \N__7534\,
            I => \N__7531\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__7531\,
            I => \uart_tx_inst.data_reg_0\
        );

    \I__1689\ : InMux
    port map (
            O => \N__7528\,
            I => \N__7515\
        );

    \I__1688\ : InMux
    port map (
            O => \N__7527\,
            I => \N__7498\
        );

    \I__1687\ : InMux
    port map (
            O => \N__7526\,
            I => \N__7498\
        );

    \I__1686\ : InMux
    port map (
            O => \N__7525\,
            I => \N__7498\
        );

    \I__1685\ : InMux
    port map (
            O => \N__7524\,
            I => \N__7498\
        );

    \I__1684\ : InMux
    port map (
            O => \N__7523\,
            I => \N__7498\
        );

    \I__1683\ : InMux
    port map (
            O => \N__7522\,
            I => \N__7498\
        );

    \I__1682\ : InMux
    port map (
            O => \N__7521\,
            I => \N__7498\
        );

    \I__1681\ : InMux
    port map (
            O => \N__7520\,
            I => \N__7498\
        );

    \I__1680\ : InMux
    port map (
            O => \N__7519\,
            I => \N__7493\
        );

    \I__1679\ : InMux
    port map (
            O => \N__7518\,
            I => \N__7493\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__7515\,
            I => \N__7490\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__7498\,
            I => \N__7487\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__7493\,
            I => \N__7478\
        );

    \I__1675\ : Span12Mux_v
    port map (
            O => \N__7490\,
            I => \N__7475\
        );

    \I__1674\ : Span4Mux_s1_h
    port map (
            O => \N__7487\,
            I => \N__7472\
        );

    \I__1673\ : InMux
    port map (
            O => \N__7486\,
            I => \N__7469\
        );

    \I__1672\ : InMux
    port map (
            O => \N__7485\,
            I => \N__7466\
        );

    \I__1671\ : InMux
    port map (
            O => \N__7484\,
            I => \N__7463\
        );

    \I__1670\ : InMux
    port map (
            O => \N__7483\,
            I => \N__7456\
        );

    \I__1669\ : InMux
    port map (
            O => \N__7482\,
            I => \N__7456\
        );

    \I__1668\ : InMux
    port map (
            O => \N__7481\,
            I => \N__7456\
        );

    \I__1667\ : Odrv4
    port map (
            O => \N__7478\,
            I => \uart_tx_inst.n7\
        );

    \I__1666\ : Odrv12
    port map (
            O => \N__7475\,
            I => \uart_tx_inst.n7\
        );

    \I__1665\ : Odrv4
    port map (
            O => \N__7472\,
            I => \uart_tx_inst.n7\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__7469\,
            I => \uart_tx_inst.n7\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__7466\,
            I => \uart_tx_inst.n7\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__7463\,
            I => \uart_tx_inst.n7\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__7456\,
            I => \uart_tx_inst.n7\
        );

    \I__1660\ : InMux
    port map (
            O => \N__7441\,
            I => \N__7438\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__7438\,
            I => \N__7433\
        );

    \I__1658\ : InMux
    port map (
            O => \N__7437\,
            I => \N__7425\
        );

    \I__1657\ : InMux
    port map (
            O => \N__7436\,
            I => \N__7425\
        );

    \I__1656\ : Span4Mux_s3_h
    port map (
            O => \N__7433\,
            I => \N__7422\
        );

    \I__1655\ : InMux
    port map (
            O => \N__7432\,
            I => \N__7419\
        );

    \I__1654\ : InMux
    port map (
            O => \N__7431\,
            I => \N__7414\
        );

    \I__1653\ : InMux
    port map (
            O => \N__7430\,
            I => \N__7414\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__7425\,
            I => \uart_tx_inst.n15\
        );

    \I__1651\ : Odrv4
    port map (
            O => \N__7422\,
            I => \uart_tx_inst.n15\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__7419\,
            I => \uart_tx_inst.n15\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__7414\,
            I => \uart_tx_inst.n15\
        );

    \I__1648\ : IoInMux
    port map (
            O => \N__7405\,
            I => \N__7402\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__7402\,
            I => \N__7399\
        );

    \I__1646\ : IoSpan4Mux
    port map (
            O => \N__7399\,
            I => \N__7396\
        );

    \I__1645\ : Span4Mux_s3_v
    port map (
            O => \N__7396\,
            I => \N__7393\
        );

    \I__1644\ : Span4Mux_v
    port map (
            O => \N__7393\,
            I => \N__7390\
        );

    \I__1643\ : Span4Mux_v
    port map (
            O => \N__7390\,
            I => \N__7387\
        );

    \I__1642\ : Odrv4
    port map (
            O => \N__7387\,
            I => txd_c
        );

    \I__1641\ : ClkMux
    port map (
            O => \N__7384\,
            I => \N__7285\
        );

    \I__1640\ : ClkMux
    port map (
            O => \N__7383\,
            I => \N__7285\
        );

    \I__1639\ : ClkMux
    port map (
            O => \N__7382\,
            I => \N__7285\
        );

    \I__1638\ : ClkMux
    port map (
            O => \N__7381\,
            I => \N__7285\
        );

    \I__1637\ : ClkMux
    port map (
            O => \N__7380\,
            I => \N__7285\
        );

    \I__1636\ : ClkMux
    port map (
            O => \N__7379\,
            I => \N__7285\
        );

    \I__1635\ : ClkMux
    port map (
            O => \N__7378\,
            I => \N__7285\
        );

    \I__1634\ : ClkMux
    port map (
            O => \N__7377\,
            I => \N__7285\
        );

    \I__1633\ : ClkMux
    port map (
            O => \N__7376\,
            I => \N__7285\
        );

    \I__1632\ : ClkMux
    port map (
            O => \N__7375\,
            I => \N__7285\
        );

    \I__1631\ : ClkMux
    port map (
            O => \N__7374\,
            I => \N__7285\
        );

    \I__1630\ : ClkMux
    port map (
            O => \N__7373\,
            I => \N__7285\
        );

    \I__1629\ : ClkMux
    port map (
            O => \N__7372\,
            I => \N__7285\
        );

    \I__1628\ : ClkMux
    port map (
            O => \N__7371\,
            I => \N__7285\
        );

    \I__1627\ : ClkMux
    port map (
            O => \N__7370\,
            I => \N__7285\
        );

    \I__1626\ : ClkMux
    port map (
            O => \N__7369\,
            I => \N__7285\
        );

    \I__1625\ : ClkMux
    port map (
            O => \N__7368\,
            I => \N__7285\
        );

    \I__1624\ : ClkMux
    port map (
            O => \N__7367\,
            I => \N__7285\
        );

    \I__1623\ : ClkMux
    port map (
            O => \N__7366\,
            I => \N__7285\
        );

    \I__1622\ : ClkMux
    port map (
            O => \N__7365\,
            I => \N__7285\
        );

    \I__1621\ : ClkMux
    port map (
            O => \N__7364\,
            I => \N__7285\
        );

    \I__1620\ : ClkMux
    port map (
            O => \N__7363\,
            I => \N__7285\
        );

    \I__1619\ : ClkMux
    port map (
            O => \N__7362\,
            I => \N__7285\
        );

    \I__1618\ : ClkMux
    port map (
            O => \N__7361\,
            I => \N__7285\
        );

    \I__1617\ : ClkMux
    port map (
            O => \N__7360\,
            I => \N__7285\
        );

    \I__1616\ : ClkMux
    port map (
            O => \N__7359\,
            I => \N__7285\
        );

    \I__1615\ : ClkMux
    port map (
            O => \N__7358\,
            I => \N__7285\
        );

    \I__1614\ : ClkMux
    port map (
            O => \N__7357\,
            I => \N__7285\
        );

    \I__1613\ : ClkMux
    port map (
            O => \N__7356\,
            I => \N__7285\
        );

    \I__1612\ : ClkMux
    port map (
            O => \N__7355\,
            I => \N__7285\
        );

    \I__1611\ : ClkMux
    port map (
            O => \N__7354\,
            I => \N__7285\
        );

    \I__1610\ : ClkMux
    port map (
            O => \N__7353\,
            I => \N__7285\
        );

    \I__1609\ : ClkMux
    port map (
            O => \N__7352\,
            I => \N__7285\
        );

    \I__1608\ : GlobalMux
    port map (
            O => \N__7285\,
            I => \N__7282\
        );

    \I__1607\ : gio2CtrlBuf
    port map (
            O => \N__7282\,
            I => clk_c
        );

    \I__1606\ : CEMux
    port map (
            O => \N__7279\,
            I => \N__7276\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__7276\,
            I => \N__7273\
        );

    \I__1604\ : Sp12to4
    port map (
            O => \N__7273\,
            I => \N__7270\
        );

    \I__1603\ : Odrv12
    port map (
            O => \N__7270\,
            I => \uart_tx_inst.n719\
        );

    \I__1602\ : SRMux
    port map (
            O => \N__7267\,
            I => \N__7259\
        );

    \I__1601\ : SRMux
    port map (
            O => \N__7266\,
            I => \N__7256\
        );

    \I__1600\ : SRMux
    port map (
            O => \N__7265\,
            I => \N__7249\
        );

    \I__1599\ : SRMux
    port map (
            O => \N__7264\,
            I => \N__7246\
        );

    \I__1598\ : CascadeMux
    port map (
            O => \N__7263\,
            I => \N__7233\
        );

    \I__1597\ : SRMux
    port map (
            O => \N__7262\,
            I => \N__7228\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__7259\,
            I => \N__7224\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__7256\,
            I => \N__7221\
        );

    \I__1594\ : InMux
    port map (
            O => \N__7255\,
            I => \N__7218\
        );

    \I__1593\ : SRMux
    port map (
            O => \N__7254\,
            I => \N__7215\
        );

    \I__1592\ : InMux
    port map (
            O => \N__7253\,
            I => \N__7212\
        );

    \I__1591\ : InMux
    port map (
            O => \N__7252\,
            I => \N__7209\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__7249\,
            I => \N__7206\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__7246\,
            I => \N__7203\
        );

    \I__1588\ : InMux
    port map (
            O => \N__7245\,
            I => \N__7200\
        );

    \I__1587\ : SRMux
    port map (
            O => \N__7244\,
            I => \N__7197\
        );

    \I__1586\ : InMux
    port map (
            O => \N__7243\,
            I => \N__7192\
        );

    \I__1585\ : InMux
    port map (
            O => \N__7242\,
            I => \N__7192\
        );

    \I__1584\ : SRMux
    port map (
            O => \N__7241\,
            I => \N__7189\
        );

    \I__1583\ : CascadeMux
    port map (
            O => \N__7240\,
            I => \N__7182\
        );

    \I__1582\ : SRMux
    port map (
            O => \N__7239\,
            I => \N__7178\
        );

    \I__1581\ : InMux
    port map (
            O => \N__7238\,
            I => \N__7172\
        );

    \I__1580\ : SRMux
    port map (
            O => \N__7237\,
            I => \N__7169\
        );

    \I__1579\ : InMux
    port map (
            O => \N__7236\,
            I => \N__7164\
        );

    \I__1578\ : InMux
    port map (
            O => \N__7233\,
            I => \N__7164\
        );

    \I__1577\ : SRMux
    port map (
            O => \N__7232\,
            I => \N__7158\
        );

    \I__1576\ : SRMux
    port map (
            O => \N__7231\,
            I => \N__7155\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__7228\,
            I => \N__7152\
        );

    \I__1574\ : SRMux
    port map (
            O => \N__7227\,
            I => \N__7149\
        );

    \I__1573\ : Span4Mux_v
    port map (
            O => \N__7224\,
            I => \N__7140\
        );

    \I__1572\ : Span4Mux_v
    port map (
            O => \N__7221\,
            I => \N__7140\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__7218\,
            I => \N__7140\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__7215\,
            I => \N__7140\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__7212\,
            I => \N__7137\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__7209\,
            I => \N__7134\
        );

    \I__1567\ : Span4Mux_v
    port map (
            O => \N__7206\,
            I => \N__7123\
        );

    \I__1566\ : Span4Mux_h
    port map (
            O => \N__7203\,
            I => \N__7123\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__7200\,
            I => \N__7123\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__7197\,
            I => \N__7123\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__7192\,
            I => \N__7118\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__7189\,
            I => \N__7118\
        );

    \I__1561\ : SRMux
    port map (
            O => \N__7188\,
            I => \N__7115\
        );

    \I__1560\ : InMux
    port map (
            O => \N__7187\,
            I => \N__7108\
        );

    \I__1559\ : InMux
    port map (
            O => \N__7186\,
            I => \N__7108\
        );

    \I__1558\ : InMux
    port map (
            O => \N__7185\,
            I => \N__7108\
        );

    \I__1557\ : InMux
    port map (
            O => \N__7182\,
            I => \N__7105\
        );

    \I__1556\ : SRMux
    port map (
            O => \N__7181\,
            I => \N__7102\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__7178\,
            I => \N__7099\
        );

    \I__1554\ : InMux
    port map (
            O => \N__7177\,
            I => \N__7096\
        );

    \I__1553\ : InMux
    port map (
            O => \N__7176\,
            I => \N__7093\
        );

    \I__1552\ : SRMux
    port map (
            O => \N__7175\,
            I => \N__7090\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__7172\,
            I => \N__7087\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__7169\,
            I => \N__7082\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__7164\,
            I => \N__7082\
        );

    \I__1548\ : SRMux
    port map (
            O => \N__7163\,
            I => \N__7079\
        );

    \I__1547\ : InMux
    port map (
            O => \N__7162\,
            I => \N__7074\
        );

    \I__1546\ : InMux
    port map (
            O => \N__7161\,
            I => \N__7074\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__7158\,
            I => \N__7069\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__7155\,
            I => \N__7066\
        );

    \I__1543\ : Span4Mux_v
    port map (
            O => \N__7152\,
            I => \N__7061\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__7149\,
            I => \N__7061\
        );

    \I__1541\ : Span4Mux_v
    port map (
            O => \N__7140\,
            I => \N__7054\
        );

    \I__1540\ : Span4Mux_h
    port map (
            O => \N__7137\,
            I => \N__7054\
        );

    \I__1539\ : Span4Mux_h
    port map (
            O => \N__7134\,
            I => \N__7054\
        );

    \I__1538\ : InMux
    port map (
            O => \N__7133\,
            I => \N__7051\
        );

    \I__1537\ : SRMux
    port map (
            O => \N__7132\,
            I => \N__7048\
        );

    \I__1536\ : Span4Mux_v
    port map (
            O => \N__7123\,
            I => \N__7043\
        );

    \I__1535\ : Span4Mux_h
    port map (
            O => \N__7118\,
            I => \N__7043\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__7115\,
            I => \N__7040\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__7108\,
            I => \N__7037\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__7105\,
            I => \N__7032\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__7102\,
            I => \N__7032\
        );

    \I__1530\ : Span4Mux_h
    port map (
            O => \N__7099\,
            I => \N__7023\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__7096\,
            I => \N__7023\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__7093\,
            I => \N__7023\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__7090\,
            I => \N__7023\
        );

    \I__1526\ : Span4Mux_v
    port map (
            O => \N__7087\,
            I => \N__7016\
        );

    \I__1525\ : Span4Mux_h
    port map (
            O => \N__7082\,
            I => \N__7016\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__7079\,
            I => \N__7016\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__7074\,
            I => \N__7013\
        );

    \I__1522\ : InMux
    port map (
            O => \N__7073\,
            I => \N__7008\
        );

    \I__1521\ : SRMux
    port map (
            O => \N__7072\,
            I => \N__7008\
        );

    \I__1520\ : Span12Mux_s8_h
    port map (
            O => \N__7069\,
            I => \N__7005\
        );

    \I__1519\ : Span12Mux_s8_h
    port map (
            O => \N__7066\,
            I => \N__7002\
        );

    \I__1518\ : IoSpan4Mux
    port map (
            O => \N__7061\,
            I => \N__6999\
        );

    \I__1517\ : Span4Mux_v
    port map (
            O => \N__7054\,
            I => \N__6992\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__7051\,
            I => \N__6992\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__7048\,
            I => \N__6992\
        );

    \I__1514\ : Span4Mux_v
    port map (
            O => \N__7043\,
            I => \N__6981\
        );

    \I__1513\ : Span4Mux_h
    port map (
            O => \N__7040\,
            I => \N__6981\
        );

    \I__1512\ : Span4Mux_h
    port map (
            O => \N__7037\,
            I => \N__6981\
        );

    \I__1511\ : Span4Mux_s3_h
    port map (
            O => \N__7032\,
            I => \N__6981\
        );

    \I__1510\ : Span4Mux_v
    port map (
            O => \N__7023\,
            I => \N__6981\
        );

    \I__1509\ : Span4Mux_v
    port map (
            O => \N__7016\,
            I => \N__6974\
        );

    \I__1508\ : Span4Mux_h
    port map (
            O => \N__7013\,
            I => \N__6974\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__7008\,
            I => \N__6974\
        );

    \I__1506\ : Odrv12
    port map (
            O => \N__7005\,
            I => rst_c
        );

    \I__1505\ : Odrv12
    port map (
            O => \N__7002\,
            I => rst_c
        );

    \I__1504\ : Odrv4
    port map (
            O => \N__6999\,
            I => rst_c
        );

    \I__1503\ : Odrv4
    port map (
            O => \N__6992\,
            I => rst_c
        );

    \I__1502\ : Odrv4
    port map (
            O => \N__6981\,
            I => rst_c
        );

    \I__1501\ : Odrv4
    port map (
            O => \N__6974\,
            I => rst_c
        );

    \I__1500\ : InMux
    port map (
            O => \N__6961\,
            I => \N__6957\
        );

    \I__1499\ : InMux
    port map (
            O => \N__6960\,
            I => \N__6954\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__6957\,
            I => \N__6951\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__6954\,
            I => \N__6948\
        );

    \I__1496\ : Span4Mux_v
    port map (
            O => \N__6951\,
            I => \N__6945\
        );

    \I__1495\ : Span4Mux_s2_v
    port map (
            O => \N__6948\,
            I => \N__6942\
        );

    \I__1494\ : Odrv4
    port map (
            O => \N__6945\,
            I => n108
        );

    \I__1493\ : Odrv4
    port map (
            O => \N__6942\,
            I => n108
        );

    \I__1492\ : InMux
    port map (
            O => \N__6937\,
            I => \bfn_12_5_0_\
        );

    \I__1491\ : InMux
    port map (
            O => \N__6934\,
            I => \N__6931\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__6931\,
            I => \N__6927\
        );

    \I__1489\ : InMux
    port map (
            O => \N__6930\,
            I => \N__6924\
        );

    \I__1488\ : Span4Mux_v
    port map (
            O => \N__6927\,
            I => \N__6921\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__6924\,
            I => \N__6918\
        );

    \I__1486\ : Span4Mux_h
    port map (
            O => \N__6921\,
            I => \N__6915\
        );

    \I__1485\ : Span4Mux_s1_v
    port map (
            O => \N__6918\,
            I => \N__6912\
        );

    \I__1484\ : Odrv4
    port map (
            O => \N__6915\,
            I => n107
        );

    \I__1483\ : Odrv4
    port map (
            O => \N__6912\,
            I => n107
        );

    \I__1482\ : InMux
    port map (
            O => \N__6907\,
            I => \uart_tx_inst.n1582\
        );

    \I__1481\ : InMux
    port map (
            O => \N__6904\,
            I => \N__6901\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__6901\,
            I => \N__6898\
        );

    \I__1479\ : Span4Mux_v
    port map (
            O => \N__6898\,
            I => \N__6894\
        );

    \I__1478\ : InMux
    port map (
            O => \N__6897\,
            I => \N__6891\
        );

    \I__1477\ : Span4Mux_h
    port map (
            O => \N__6894\,
            I => \N__6888\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__6891\,
            I => \N__6885\
        );

    \I__1475\ : Odrv4
    port map (
            O => \N__6888\,
            I => n106
        );

    \I__1474\ : Odrv12
    port map (
            O => \N__6885\,
            I => n106
        );

    \I__1473\ : CascadeMux
    port map (
            O => \N__6880\,
            I => \uart_tx_inst.n865_cascade_\
        );

    \I__1472\ : CascadeMux
    port map (
            O => \N__6877\,
            I => \N__6874\
        );

    \I__1471\ : InMux
    port map (
            O => \N__6874\,
            I => \N__6870\
        );

    \I__1470\ : InMux
    port map (
            O => \N__6873\,
            I => \N__6867\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__6870\,
            I => \uart_tx_inst.prescale_reg_4\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__6867\,
            I => \uart_tx_inst.prescale_reg_4\
        );

    \I__1467\ : CascadeMux
    port map (
            O => \N__6862\,
            I => \N__6859\
        );

    \I__1466\ : InMux
    port map (
            O => \N__6859\,
            I => \N__6856\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__6856\,
            I => \uart_tx_inst.n31\
        );

    \I__1464\ : CascadeMux
    port map (
            O => \N__6853\,
            I => \uart_tx_inst.n870_cascade_\
        );

    \I__1463\ : InMux
    port map (
            O => \N__6850\,
            I => \N__6846\
        );

    \I__1462\ : InMux
    port map (
            O => \N__6849\,
            I => \N__6843\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__6846\,
            I => \uart_tx_inst.prescale_reg_5\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__6843\,
            I => \uart_tx_inst.prescale_reg_5\
        );

    \I__1459\ : InMux
    port map (
            O => \N__6838\,
            I => \N__6827\
        );

    \I__1458\ : InMux
    port map (
            O => \N__6837\,
            I => \N__6827\
        );

    \I__1457\ : InMux
    port map (
            O => \N__6836\,
            I => \N__6824\
        );

    \I__1456\ : InMux
    port map (
            O => \N__6835\,
            I => \N__6821\
        );

    \I__1455\ : InMux
    port map (
            O => \N__6834\,
            I => \N__6816\
        );

    \I__1454\ : InMux
    port map (
            O => \N__6833\,
            I => \N__6816\
        );

    \I__1453\ : CascadeMux
    port map (
            O => \N__6832\,
            I => \N__6813\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__6827\,
            I => \N__6799\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__6824\,
            I => \N__6799\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__6821\,
            I => \N__6794\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__6816\,
            I => \N__6794\
        );

    \I__1448\ : InMux
    port map (
            O => \N__6813\,
            I => \N__6787\
        );

    \I__1447\ : InMux
    port map (
            O => \N__6812\,
            I => \N__6787\
        );

    \I__1446\ : InMux
    port map (
            O => \N__6811\,
            I => \N__6787\
        );

    \I__1445\ : InMux
    port map (
            O => \N__6810\,
            I => \N__6778\
        );

    \I__1444\ : InMux
    port map (
            O => \N__6809\,
            I => \N__6778\
        );

    \I__1443\ : InMux
    port map (
            O => \N__6808\,
            I => \N__6778\
        );

    \I__1442\ : InMux
    port map (
            O => \N__6807\,
            I => \N__6778\
        );

    \I__1441\ : InMux
    port map (
            O => \N__6806\,
            I => \N__6767\
        );

    \I__1440\ : InMux
    port map (
            O => \N__6805\,
            I => \N__6767\
        );

    \I__1439\ : InMux
    port map (
            O => \N__6804\,
            I => \N__6767\
        );

    \I__1438\ : Span4Mux_s3_h
    port map (
            O => \N__6799\,
            I => \N__6764\
        );

    \I__1437\ : Span4Mux_v
    port map (
            O => \N__6794\,
            I => \N__6761\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__6787\,
            I => \N__6756\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__6778\,
            I => \N__6756\
        );

    \I__1434\ : InMux
    port map (
            O => \N__6777\,
            I => \N__6747\
        );

    \I__1433\ : InMux
    port map (
            O => \N__6776\,
            I => \N__6747\
        );

    \I__1432\ : InMux
    port map (
            O => \N__6775\,
            I => \N__6747\
        );

    \I__1431\ : InMux
    port map (
            O => \N__6774\,
            I => \N__6747\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__6767\,
            I => \uart_tx_inst.n485\
        );

    \I__1429\ : Odrv4
    port map (
            O => \N__6764\,
            I => \uart_tx_inst.n485\
        );

    \I__1428\ : Odrv4
    port map (
            O => \N__6761\,
            I => \uart_tx_inst.n485\
        );

    \I__1427\ : Odrv12
    port map (
            O => \N__6756\,
            I => \uart_tx_inst.n485\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__6747\,
            I => \uart_tx_inst.n485\
        );

    \I__1425\ : InMux
    port map (
            O => \N__6736\,
            I => \N__6733\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__6733\,
            I => \N__6730\
        );

    \I__1423\ : Odrv4
    port map (
            O => \N__6730\,
            I => \uart_tx_inst.n28\
        );

    \I__1422\ : InMux
    port map (
            O => \N__6727\,
            I => \N__6714\
        );

    \I__1421\ : InMux
    port map (
            O => \N__6726\,
            I => \N__6714\
        );

    \I__1420\ : InMux
    port map (
            O => \N__6725\,
            I => \N__6714\
        );

    \I__1419\ : InMux
    port map (
            O => \N__6724\,
            I => \N__6700\
        );

    \I__1418\ : InMux
    port map (
            O => \N__6723\,
            I => \N__6700\
        );

    \I__1417\ : InMux
    port map (
            O => \N__6722\,
            I => \N__6700\
        );

    \I__1416\ : InMux
    port map (
            O => \N__6721\,
            I => \N__6693\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__6714\,
            I => \N__6686\
        );

    \I__1414\ : InMux
    port map (
            O => \N__6713\,
            I => \N__6677\
        );

    \I__1413\ : InMux
    port map (
            O => \N__6712\,
            I => \N__6677\
        );

    \I__1412\ : InMux
    port map (
            O => \N__6711\,
            I => \N__6677\
        );

    \I__1411\ : InMux
    port map (
            O => \N__6710\,
            I => \N__6677\
        );

    \I__1410\ : InMux
    port map (
            O => \N__6709\,
            I => \N__6670\
        );

    \I__1409\ : InMux
    port map (
            O => \N__6708\,
            I => \N__6670\
        );

    \I__1408\ : InMux
    port map (
            O => \N__6707\,
            I => \N__6670\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__6700\,
            I => \N__6664\
        );

    \I__1406\ : InMux
    port map (
            O => \N__6699\,
            I => \N__6655\
        );

    \I__1405\ : InMux
    port map (
            O => \N__6698\,
            I => \N__6655\
        );

    \I__1404\ : InMux
    port map (
            O => \N__6697\,
            I => \N__6655\
        );

    \I__1403\ : InMux
    port map (
            O => \N__6696\,
            I => \N__6655\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__6693\,
            I => \N__6652\
        );

    \I__1401\ : InMux
    port map (
            O => \N__6692\,
            I => \N__6643\
        );

    \I__1400\ : InMux
    port map (
            O => \N__6691\,
            I => \N__6643\
        );

    \I__1399\ : InMux
    port map (
            O => \N__6690\,
            I => \N__6643\
        );

    \I__1398\ : InMux
    port map (
            O => \N__6689\,
            I => \N__6643\
        );

    \I__1397\ : Span4Mux_s0_h
    port map (
            O => \N__6686\,
            I => \N__6638\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__6677\,
            I => \N__6638\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__6670\,
            I => \N__6635\
        );

    \I__1394\ : InMux
    port map (
            O => \N__6669\,
            I => \N__6632\
        );

    \I__1393\ : InMux
    port map (
            O => \N__6668\,
            I => \N__6629\
        );

    \I__1392\ : InMux
    port map (
            O => \N__6667\,
            I => \N__6626\
        );

    \I__1391\ : Odrv4
    port map (
            O => \N__6664\,
            I => \input_axis_tready_N_72\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__6655\,
            I => \input_axis_tready_N_72\
        );

    \I__1389\ : Odrv4
    port map (
            O => \N__6652\,
            I => \input_axis_tready_N_72\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__6643\,
            I => \input_axis_tready_N_72\
        );

    \I__1387\ : Odrv4
    port map (
            O => \N__6638\,
            I => \input_axis_tready_N_72\
        );

    \I__1386\ : Odrv4
    port map (
            O => \N__6635\,
            I => \input_axis_tready_N_72\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__6632\,
            I => \input_axis_tready_N_72\
        );

    \I__1384\ : LocalMux
    port map (
            O => \N__6629\,
            I => \input_axis_tready_N_72\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__6626\,
            I => \input_axis_tready_N_72\
        );

    \I__1382\ : CascadeMux
    port map (
            O => \N__6607\,
            I => \uart_tx_inst.n885_cascade_\
        );

    \I__1381\ : InMux
    port map (
            O => \N__6604\,
            I => \N__6598\
        );

    \I__1380\ : InMux
    port map (
            O => \N__6603\,
            I => \N__6598\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__6598\,
            I => \N__6589\
        );

    \I__1378\ : InMux
    port map (
            O => \N__6597\,
            I => \N__6586\
        );

    \I__1377\ : InMux
    port map (
            O => \N__6596\,
            I => \N__6577\
        );

    \I__1376\ : InMux
    port map (
            O => \N__6595\,
            I => \N__6577\
        );

    \I__1375\ : InMux
    port map (
            O => \N__6594\,
            I => \N__6577\
        );

    \I__1374\ : InMux
    port map (
            O => \N__6593\,
            I => \N__6577\
        );

    \I__1373\ : CascadeMux
    port map (
            O => \N__6592\,
            I => \N__6563\
        );

    \I__1372\ : Span4Mux_s1_v
    port map (
            O => \N__6589\,
            I => \N__6560\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__6586\,
            I => \N__6555\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__6577\,
            I => \N__6555\
        );

    \I__1369\ : InMux
    port map (
            O => \N__6576\,
            I => \N__6551\
        );

    \I__1368\ : InMux
    port map (
            O => \N__6575\,
            I => \N__6544\
        );

    \I__1367\ : InMux
    port map (
            O => \N__6574\,
            I => \N__6544\
        );

    \I__1366\ : InMux
    port map (
            O => \N__6573\,
            I => \N__6544\
        );

    \I__1365\ : InMux
    port map (
            O => \N__6572\,
            I => \N__6539\
        );

    \I__1364\ : InMux
    port map (
            O => \N__6571\,
            I => \N__6539\
        );

    \I__1363\ : InMux
    port map (
            O => \N__6570\,
            I => \N__6536\
        );

    \I__1362\ : InMux
    port map (
            O => \N__6569\,
            I => \N__6533\
        );

    \I__1361\ : InMux
    port map (
            O => \N__6568\,
            I => \N__6524\
        );

    \I__1360\ : InMux
    port map (
            O => \N__6567\,
            I => \N__6524\
        );

    \I__1359\ : InMux
    port map (
            O => \N__6566\,
            I => \N__6524\
        );

    \I__1358\ : InMux
    port map (
            O => \N__6563\,
            I => \N__6524\
        );

    \I__1357\ : Span4Mux_s0_h
    port map (
            O => \N__6560\,
            I => \N__6519\
        );

    \I__1356\ : Span4Mux_s1_v
    port map (
            O => \N__6555\,
            I => \N__6519\
        );

    \I__1355\ : InMux
    port map (
            O => \N__6554\,
            I => \N__6516\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__6551\,
            I => \uart_tx_inst.n165\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__6544\,
            I => \uart_tx_inst.n165\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__6539\,
            I => \uart_tx_inst.n165\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__6536\,
            I => \uart_tx_inst.n165\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__6533\,
            I => \uart_tx_inst.n165\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__6524\,
            I => \uart_tx_inst.n165\
        );

    \I__1348\ : Odrv4
    port map (
            O => \N__6519\,
            I => \uart_tx_inst.n165\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__6516\,
            I => \uart_tx_inst.n165\
        );

    \I__1346\ : InMux
    port map (
            O => \N__6499\,
            I => \N__6495\
        );

    \I__1345\ : CascadeMux
    port map (
            O => \N__6498\,
            I => \N__6492\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__6495\,
            I => \N__6489\
        );

    \I__1343\ : InMux
    port map (
            O => \N__6492\,
            I => \N__6486\
        );

    \I__1342\ : Odrv4
    port map (
            O => \N__6489\,
            I => \uart_tx_inst.prescale_reg_8\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__6486\,
            I => \uart_tx_inst.prescale_reg_8\
        );

    \I__1340\ : CEMux
    port map (
            O => \N__6481\,
            I => \N__6478\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__6478\,
            I => \N__6472\
        );

    \I__1338\ : CEMux
    port map (
            O => \N__6477\,
            I => \N__6469\
        );

    \I__1337\ : CEMux
    port map (
            O => \N__6476\,
            I => \N__6466\
        );

    \I__1336\ : CEMux
    port map (
            O => \N__6475\,
            I => \N__6461\
        );

    \I__1335\ : Span4Mux_v
    port map (
            O => \N__6472\,
            I => \N__6454\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__6469\,
            I => \N__6454\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__6466\,
            I => \N__6454\
        );

    \I__1332\ : CEMux
    port map (
            O => \N__6465\,
            I => \N__6451\
        );

    \I__1331\ : CEMux
    port map (
            O => \N__6464\,
            I => \N__6448\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__6461\,
            I => \N__6445\
        );

    \I__1329\ : Span4Mux_h
    port map (
            O => \N__6454\,
            I => \N__6442\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__6451\,
            I => \N__6439\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__6448\,
            I => \N__6436\
        );

    \I__1326\ : Span4Mux_s0_v
    port map (
            O => \N__6445\,
            I => \N__6431\
        );

    \I__1325\ : Span4Mux_s0_h
    port map (
            O => \N__6442\,
            I => \N__6431\
        );

    \I__1324\ : Odrv12
    port map (
            O => \N__6439\,
            I => \uart_tx_inst.n873\
        );

    \I__1323\ : Odrv4
    port map (
            O => \N__6436\,
            I => \uart_tx_inst.n873\
        );

    \I__1322\ : Odrv4
    port map (
            O => \N__6431\,
            I => \uart_tx_inst.n873\
        );

    \I__1321\ : InMux
    port map (
            O => \N__6424\,
            I => \N__6421\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__6421\,
            I => \uart_tx_inst.data_reg_1\
        );

    \I__1319\ : InMux
    port map (
            O => \N__6418\,
            I => \N__6415\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__6415\,
            I => \uart_tx_inst.data_reg_2\
        );

    \I__1317\ : InMux
    port map (
            O => \N__6412\,
            I => \N__6409\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__6409\,
            I => \N__6406\
        );

    \I__1315\ : Span4Mux_v
    port map (
            O => \N__6406\,
            I => \N__6403\
        );

    \I__1314\ : Odrv4
    port map (
            O => \N__6403\,
            I => \uart_rx_inst.n317\
        );

    \I__1313\ : InMux
    port map (
            O => \N__6400\,
            I => \uart_rx_inst.n1540\
        );

    \I__1312\ : InMux
    port map (
            O => \N__6397\,
            I => \N__6394\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__6394\,
            I => \N__6391\
        );

    \I__1310\ : Span4Mux_h
    port map (
            O => \N__6391\,
            I => \N__6388\
        );

    \I__1309\ : Odrv4
    port map (
            O => \N__6388\,
            I => \uart_rx_inst.n316\
        );

    \I__1308\ : InMux
    port map (
            O => \N__6385\,
            I => \uart_rx_inst.n1541\
        );

    \I__1307\ : InMux
    port map (
            O => \N__6382\,
            I => \N__6379\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__6379\,
            I => \N__6376\
        );

    \I__1305\ : Span4Mux_v
    port map (
            O => \N__6376\,
            I => \N__6373\
        );

    \I__1304\ : Odrv4
    port map (
            O => \N__6373\,
            I => \uart_rx_inst.n315\
        );

    \I__1303\ : InMux
    port map (
            O => \N__6370\,
            I => \uart_rx_inst.n1542\
        );

    \I__1302\ : InMux
    port map (
            O => \N__6367\,
            I => \N__6364\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__6364\,
            I => \N__6361\
        );

    \I__1300\ : Span4Mux_h
    port map (
            O => \N__6361\,
            I => \N__6358\
        );

    \I__1299\ : Odrv4
    port map (
            O => \N__6358\,
            I => \uart_rx_inst.n314\
        );

    \I__1298\ : InMux
    port map (
            O => \N__6355\,
            I => \uart_rx_inst.n1543\
        );

    \I__1297\ : InMux
    port map (
            O => \N__6352\,
            I => \N__6349\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__6349\,
            I => \N__6346\
        );

    \I__1295\ : Span4Mux_v
    port map (
            O => \N__6346\,
            I => \N__6343\
        );

    \I__1294\ : Odrv4
    port map (
            O => \N__6343\,
            I => \uart_rx_inst.n313\
        );

    \I__1293\ : InMux
    port map (
            O => \N__6340\,
            I => \uart_rx_inst.n1544\
        );

    \I__1292\ : InMux
    port map (
            O => \N__6337\,
            I => \bfn_11_7_0_\
        );

    \I__1291\ : InMux
    port map (
            O => \N__6334\,
            I => \N__6331\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__6331\,
            I => \N__6328\
        );

    \I__1289\ : Span4Mux_v
    port map (
            O => \N__6328\,
            I => \N__6325\
        );

    \I__1288\ : Odrv4
    port map (
            O => \N__6325\,
            I => \uart_rx_inst.n312\
        );

    \I__1287\ : InMux
    port map (
            O => \N__6322\,
            I => \N__6315\
        );

    \I__1286\ : InMux
    port map (
            O => \N__6321\,
            I => \N__6315\
        );

    \I__1285\ : InMux
    port map (
            O => \N__6320\,
            I => \N__6308\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__6315\,
            I => \N__6305\
        );

    \I__1283\ : InMux
    port map (
            O => \N__6314\,
            I => \N__6289\
        );

    \I__1282\ : InMux
    port map (
            O => \N__6313\,
            I => \N__6282\
        );

    \I__1281\ : InMux
    port map (
            O => \N__6312\,
            I => \N__6282\
        );

    \I__1280\ : InMux
    port map (
            O => \N__6311\,
            I => \N__6279\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__6308\,
            I => \N__6276\
        );

    \I__1278\ : Span4Mux_v
    port map (
            O => \N__6305\,
            I => \N__6273\
        );

    \I__1277\ : InMux
    port map (
            O => \N__6304\,
            I => \N__6262\
        );

    \I__1276\ : InMux
    port map (
            O => \N__6303\,
            I => \N__6262\
        );

    \I__1275\ : InMux
    port map (
            O => \N__6302\,
            I => \N__6262\
        );

    \I__1274\ : InMux
    port map (
            O => \N__6301\,
            I => \N__6262\
        );

    \I__1273\ : InMux
    port map (
            O => \N__6300\,
            I => \N__6262\
        );

    \I__1272\ : InMux
    port map (
            O => \N__6299\,
            I => \N__6245\
        );

    \I__1271\ : InMux
    port map (
            O => \N__6298\,
            I => \N__6245\
        );

    \I__1270\ : InMux
    port map (
            O => \N__6297\,
            I => \N__6245\
        );

    \I__1269\ : InMux
    port map (
            O => \N__6296\,
            I => \N__6245\
        );

    \I__1268\ : InMux
    port map (
            O => \N__6295\,
            I => \N__6245\
        );

    \I__1267\ : InMux
    port map (
            O => \N__6294\,
            I => \N__6245\
        );

    \I__1266\ : InMux
    port map (
            O => \N__6293\,
            I => \N__6245\
        );

    \I__1265\ : InMux
    port map (
            O => \N__6292\,
            I => \N__6245\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__6289\,
            I => \N__6242\
        );

    \I__1263\ : InMux
    port map (
            O => \N__6288\,
            I => \N__6237\
        );

    \I__1262\ : InMux
    port map (
            O => \N__6287\,
            I => \N__6237\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__6282\,
            I => \uart_rx_inst.n232\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__6279\,
            I => \uart_rx_inst.n232\
        );

    \I__1259\ : Odrv4
    port map (
            O => \N__6276\,
            I => \uart_rx_inst.n232\
        );

    \I__1258\ : Odrv4
    port map (
            O => \N__6273\,
            I => \uart_rx_inst.n232\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__6262\,
            I => \uart_rx_inst.n232\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__6245\,
            I => \uart_rx_inst.n232\
        );

    \I__1255\ : Odrv4
    port map (
            O => \N__6242\,
            I => \uart_rx_inst.n232\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__6237\,
            I => \uart_rx_inst.n232\
        );

    \I__1253\ : InMux
    port map (
            O => \N__6220\,
            I => \N__6217\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__6217\,
            I => \N__6214\
        );

    \I__1251\ : Span4Mux_h
    port map (
            O => \N__6214\,
            I => \N__6211\
        );

    \I__1250\ : Odrv4
    port map (
            O => \N__6211\,
            I => \uart_rx_inst.n1746\
        );

    \I__1249\ : InMux
    port map (
            O => \N__6208\,
            I => \N__6204\
        );

    \I__1248\ : InMux
    port map (
            O => \N__6207\,
            I => \N__6201\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__6204\,
            I => \uart_tx_inst.prescale_reg_0\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__6201\,
            I => \uart_tx_inst.prescale_reg_0\
        );

    \I__1245\ : InMux
    port map (
            O => \N__6196\,
            I => \N__6193\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__6193\,
            I => \N__6190\
        );

    \I__1243\ : Odrv12
    port map (
            O => \N__6190\,
            I => \uart_tx_inst.n32_adj_197\
        );

    \I__1242\ : InMux
    port map (
            O => \N__6187\,
            I => \N__6184\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__6184\,
            I => \uart_tx_inst.n32\
        );

    \I__1240\ : InMux
    port map (
            O => \N__6181\,
            I => \N__6178\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__6178\,
            I => \N__6175\
        );

    \I__1238\ : Odrv12
    port map (
            O => \N__6175\,
            I => \uart_rx_inst.n325\
        );

    \I__1237\ : InMux
    port map (
            O => \N__6172\,
            I => \uart_rx_inst.n1532\
        );

    \I__1236\ : CascadeMux
    port map (
            O => \N__6169\,
            I => \N__6166\
        );

    \I__1235\ : InMux
    port map (
            O => \N__6166\,
            I => \N__6163\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__6163\,
            I => \N__6160\
        );

    \I__1233\ : Odrv4
    port map (
            O => \N__6160\,
            I => \uart_rx_inst.n324\
        );

    \I__1232\ : InMux
    port map (
            O => \N__6157\,
            I => \uart_rx_inst.n1533\
        );

    \I__1231\ : InMux
    port map (
            O => \N__6154\,
            I => \N__6151\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__6151\,
            I => \N__6148\
        );

    \I__1229\ : Odrv4
    port map (
            O => \N__6148\,
            I => \uart_rx_inst.n323\
        );

    \I__1228\ : InMux
    port map (
            O => \N__6145\,
            I => \uart_rx_inst.n1534\
        );

    \I__1227\ : InMux
    port map (
            O => \N__6142\,
            I => \N__6139\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__6139\,
            I => \N__6136\
        );

    \I__1225\ : Span4Mux_h
    port map (
            O => \N__6136\,
            I => \N__6133\
        );

    \I__1224\ : Odrv4
    port map (
            O => \N__6133\,
            I => \uart_rx_inst.n322\
        );

    \I__1223\ : InMux
    port map (
            O => \N__6130\,
            I => \uart_rx_inst.n1535\
        );

    \I__1222\ : InMux
    port map (
            O => \N__6127\,
            I => \N__6124\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__6124\,
            I => \N__6121\
        );

    \I__1220\ : Odrv4
    port map (
            O => \N__6121\,
            I => \uart_rx_inst.n321\
        );

    \I__1219\ : InMux
    port map (
            O => \N__6118\,
            I => \uart_rx_inst.n1536\
        );

    \I__1218\ : InMux
    port map (
            O => \N__6115\,
            I => \N__6112\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__6112\,
            I => \N__6109\
        );

    \I__1216\ : Span4Mux_v
    port map (
            O => \N__6109\,
            I => \N__6106\
        );

    \I__1215\ : Odrv4
    port map (
            O => \N__6106\,
            I => \uart_rx_inst.n320\
        );

    \I__1214\ : InMux
    port map (
            O => \N__6103\,
            I => \bfn_11_6_0_\
        );

    \I__1213\ : InMux
    port map (
            O => \N__6100\,
            I => \N__6097\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__6097\,
            I => \N__6094\
        );

    \I__1211\ : Span4Mux_v
    port map (
            O => \N__6094\,
            I => \N__6091\
        );

    \I__1210\ : Odrv4
    port map (
            O => \N__6091\,
            I => \uart_rx_inst.n319\
        );

    \I__1209\ : InMux
    port map (
            O => \N__6088\,
            I => \uart_rx_inst.n1538\
        );

    \I__1208\ : InMux
    port map (
            O => \N__6085\,
            I => \N__6082\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__6082\,
            I => \N__6079\
        );

    \I__1206\ : Span4Mux_h
    port map (
            O => \N__6079\,
            I => \N__6076\
        );

    \I__1205\ : Odrv4
    port map (
            O => \N__6076\,
            I => \uart_rx_inst.n318\
        );

    \I__1204\ : InMux
    port map (
            O => \N__6073\,
            I => \uart_rx_inst.n1539\
        );

    \I__1203\ : InMux
    port map (
            O => \N__6070\,
            I => \N__6067\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__6067\,
            I => \N__6064\
        );

    \I__1201\ : Span4Mux_s2_h
    port map (
            O => \N__6064\,
            I => \N__6060\
        );

    \I__1200\ : InMux
    port map (
            O => \N__6063\,
            I => \N__6057\
        );

    \I__1199\ : Odrv4
    port map (
            O => \N__6060\,
            I => \uart_tx_inst.prescale_reg_14\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__6057\,
            I => \uart_tx_inst.prescale_reg_14\
        );

    \I__1197\ : InMux
    port map (
            O => \N__6052\,
            I => \N__6049\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__6049\,
            I => \N__6046\
        );

    \I__1195\ : Span4Mux_s2_v
    port map (
            O => \N__6046\,
            I => \N__6043\
        );

    \I__1194\ : Odrv4
    port map (
            O => \N__6043\,
            I => \uart_tx_inst.n22\
        );

    \I__1193\ : InMux
    port map (
            O => \N__6040\,
            I => \uart_tx_inst.n1559\
        );

    \I__1192\ : CascadeMux
    port map (
            O => \N__6037\,
            I => \N__6034\
        );

    \I__1191\ : InMux
    port map (
            O => \N__6034\,
            I => \N__6031\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__6031\,
            I => \N__6028\
        );

    \I__1189\ : Span4Mux_v
    port map (
            O => \N__6028\,
            I => \N__6024\
        );

    \I__1188\ : InMux
    port map (
            O => \N__6027\,
            I => \N__6021\
        );

    \I__1187\ : Odrv4
    port map (
            O => \N__6024\,
            I => \uart_tx_inst.prescale_reg_15\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__6021\,
            I => \uart_tx_inst.prescale_reg_15\
        );

    \I__1185\ : InMux
    port map (
            O => \N__6016\,
            I => \N__6013\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__6013\,
            I => \N__6010\
        );

    \I__1183\ : Span4Mux_s2_v
    port map (
            O => \N__6010\,
            I => \N__6007\
        );

    \I__1182\ : Odrv4
    port map (
            O => \N__6007\,
            I => \uart_tx_inst.n21\
        );

    \I__1181\ : InMux
    port map (
            O => \N__6004\,
            I => \uart_tx_inst.n1560\
        );

    \I__1180\ : InMux
    port map (
            O => \N__6001\,
            I => \N__5997\
        );

    \I__1179\ : CascadeMux
    port map (
            O => \N__6000\,
            I => \N__5994\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__5997\,
            I => \N__5991\
        );

    \I__1177\ : InMux
    port map (
            O => \N__5994\,
            I => \N__5988\
        );

    \I__1176\ : Span4Mux_s2_h
    port map (
            O => \N__5991\,
            I => \N__5985\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__5988\,
            I => \N__5982\
        );

    \I__1174\ : Odrv4
    port map (
            O => \N__5985\,
            I => \uart_tx_inst.prescale_reg_16\
        );

    \I__1173\ : Odrv4
    port map (
            O => \N__5982\,
            I => \uart_tx_inst.prescale_reg_16\
        );

    \I__1172\ : InMux
    port map (
            O => \N__5977\,
            I => \N__5974\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__5974\,
            I => \N__5971\
        );

    \I__1170\ : Odrv4
    port map (
            O => \N__5971\,
            I => \uart_tx_inst.n20\
        );

    \I__1169\ : InMux
    port map (
            O => \N__5968\,
            I => \bfn_11_4_0_\
        );

    \I__1168\ : CascadeMux
    port map (
            O => \N__5965\,
            I => \N__5962\
        );

    \I__1167\ : InMux
    port map (
            O => \N__5962\,
            I => \N__5959\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__5959\,
            I => \N__5956\
        );

    \I__1165\ : Span4Mux_s2_h
    port map (
            O => \N__5956\,
            I => \N__5952\
        );

    \I__1164\ : InMux
    port map (
            O => \N__5955\,
            I => \N__5949\
        );

    \I__1163\ : Odrv4
    port map (
            O => \N__5952\,
            I => \uart_tx_inst.prescale_reg_17\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__5949\,
            I => \uart_tx_inst.prescale_reg_17\
        );

    \I__1161\ : InMux
    port map (
            O => \N__5944\,
            I => \N__5941\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__5941\,
            I => \N__5938\
        );

    \I__1159\ : Span4Mux_h
    port map (
            O => \N__5938\,
            I => \N__5935\
        );

    \I__1158\ : Odrv4
    port map (
            O => \N__5935\,
            I => \uart_tx_inst.n19\
        );

    \I__1157\ : InMux
    port map (
            O => \N__5932\,
            I => \uart_tx_inst.n1562\
        );

    \I__1156\ : InMux
    port map (
            O => \N__5929\,
            I => \N__5925\
        );

    \I__1155\ : CascadeMux
    port map (
            O => \N__5928\,
            I => \N__5922\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__5925\,
            I => \N__5919\
        );

    \I__1153\ : InMux
    port map (
            O => \N__5922\,
            I => \N__5916\
        );

    \I__1152\ : Span4Mux_v
    port map (
            O => \N__5919\,
            I => \N__5913\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__5916\,
            I => \N__5910\
        );

    \I__1150\ : Odrv4
    port map (
            O => \N__5913\,
            I => \uart_tx_inst.prescale_reg_18\
        );

    \I__1149\ : Odrv4
    port map (
            O => \N__5910\,
            I => \uart_tx_inst.prescale_reg_18\
        );

    \I__1148\ : InMux
    port map (
            O => \N__5905\,
            I => \uart_tx_inst.n1563\
        );

    \I__1147\ : InMux
    port map (
            O => \N__5902\,
            I => \N__5899\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__5899\,
            I => \N__5896\
        );

    \I__1145\ : Odrv4
    port map (
            O => \N__5896\,
            I => \uart_tx_inst.n18\
        );

    \I__1144\ : InMux
    port map (
            O => \N__5893\,
            I => \N__5890\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__5890\,
            I => \N__5887\
        );

    \I__1142\ : Span4Mux_h
    port map (
            O => \N__5887\,
            I => \N__5884\
        );

    \I__1141\ : Odrv4
    port map (
            O => \N__5884\,
            I => \uart_rx_inst.n328\
        );

    \I__1140\ : InMux
    port map (
            O => \N__5881\,
            I => \bfn_11_5_0_\
        );

    \I__1139\ : InMux
    port map (
            O => \N__5878\,
            I => \N__5875\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__5875\,
            I => \N__5872\
        );

    \I__1137\ : Odrv12
    port map (
            O => \N__5872\,
            I => \uart_rx_inst.n327\
        );

    \I__1136\ : InMux
    port map (
            O => \N__5869\,
            I => \uart_rx_inst.n1530\
        );

    \I__1135\ : InMux
    port map (
            O => \N__5866\,
            I => \N__5863\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__5863\,
            I => \N__5860\
        );

    \I__1133\ : Odrv12
    port map (
            O => \N__5860\,
            I => \uart_rx_inst.n326\
        );

    \I__1132\ : InMux
    port map (
            O => \N__5857\,
            I => \uart_rx_inst.n1531\
        );

    \I__1131\ : CascadeMux
    port map (
            O => \N__5854\,
            I => \N__5851\
        );

    \I__1130\ : InMux
    port map (
            O => \N__5851\,
            I => \N__5847\
        );

    \I__1129\ : InMux
    port map (
            O => \N__5850\,
            I => \N__5844\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__5847\,
            I => \N__5841\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__5844\,
            I => \uart_tx_inst.prescale_reg_6\
        );

    \I__1126\ : Odrv4
    port map (
            O => \N__5841\,
            I => \uart_tx_inst.prescale_reg_6\
        );

    \I__1125\ : InMux
    port map (
            O => \N__5836\,
            I => \N__5833\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__5833\,
            I => \N__5830\
        );

    \I__1123\ : Odrv12
    port map (
            O => \N__5830\,
            I => \uart_tx_inst.n30\
        );

    \I__1122\ : InMux
    port map (
            O => \N__5827\,
            I => \uart_tx_inst.n1551\
        );

    \I__1121\ : InMux
    port map (
            O => \N__5824\,
            I => \N__5820\
        );

    \I__1120\ : InMux
    port map (
            O => \N__5823\,
            I => \N__5817\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__5820\,
            I => \N__5814\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__5817\,
            I => \uart_tx_inst.prescale_reg_7\
        );

    \I__1117\ : Odrv4
    port map (
            O => \N__5814\,
            I => \uart_tx_inst.prescale_reg_7\
        );

    \I__1116\ : InMux
    port map (
            O => \N__5809\,
            I => \N__5806\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__5806\,
            I => \N__5803\
        );

    \I__1114\ : Odrv4
    port map (
            O => \N__5803\,
            I => \uart_tx_inst.n29\
        );

    \I__1113\ : InMux
    port map (
            O => \N__5800\,
            I => \uart_tx_inst.n1552\
        );

    \I__1112\ : InMux
    port map (
            O => \N__5797\,
            I => \bfn_11_3_0_\
        );

    \I__1111\ : CascadeMux
    port map (
            O => \N__5794\,
            I => \N__5791\
        );

    \I__1110\ : InMux
    port map (
            O => \N__5791\,
            I => \N__5787\
        );

    \I__1109\ : CascadeMux
    port map (
            O => \N__5790\,
            I => \N__5784\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__5787\,
            I => \N__5781\
        );

    \I__1107\ : InMux
    port map (
            O => \N__5784\,
            I => \N__5778\
        );

    \I__1106\ : Odrv4
    port map (
            O => \N__5781\,
            I => \uart_tx_inst.prescale_reg_9\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__5778\,
            I => \uart_tx_inst.prescale_reg_9\
        );

    \I__1104\ : InMux
    port map (
            O => \N__5773\,
            I => \N__5770\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__5770\,
            I => \N__5767\
        );

    \I__1102\ : Odrv4
    port map (
            O => \N__5767\,
            I => \uart_tx_inst.n27\
        );

    \I__1101\ : InMux
    port map (
            O => \N__5764\,
            I => \uart_tx_inst.n1554\
        );

    \I__1100\ : InMux
    port map (
            O => \N__5761\,
            I => \N__5758\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__5758\,
            I => \N__5755\
        );

    \I__1098\ : Span4Mux_s2_h
    port map (
            O => \N__5755\,
            I => \N__5751\
        );

    \I__1097\ : InMux
    port map (
            O => \N__5754\,
            I => \N__5748\
        );

    \I__1096\ : Odrv4
    port map (
            O => \N__5751\,
            I => \uart_tx_inst.prescale_reg_10\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__5748\,
            I => \uart_tx_inst.prescale_reg_10\
        );

    \I__1094\ : InMux
    port map (
            O => \N__5743\,
            I => \N__5740\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__5740\,
            I => \N__5737\
        );

    \I__1092\ : Span4Mux_s2_v
    port map (
            O => \N__5737\,
            I => \N__5734\
        );

    \I__1091\ : Odrv4
    port map (
            O => \N__5734\,
            I => \uart_tx_inst.n26\
        );

    \I__1090\ : InMux
    port map (
            O => \N__5731\,
            I => \uart_tx_inst.n1555\
        );

    \I__1089\ : CascadeMux
    port map (
            O => \N__5728\,
            I => \N__5725\
        );

    \I__1088\ : InMux
    port map (
            O => \N__5725\,
            I => \N__5721\
        );

    \I__1087\ : InMux
    port map (
            O => \N__5724\,
            I => \N__5718\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__5721\,
            I => \N__5715\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__5718\,
            I => \N__5712\
        );

    \I__1084\ : Odrv4
    port map (
            O => \N__5715\,
            I => \uart_tx_inst.prescale_reg_11\
        );

    \I__1083\ : Odrv4
    port map (
            O => \N__5712\,
            I => \uart_tx_inst.prescale_reg_11\
        );

    \I__1082\ : InMux
    port map (
            O => \N__5707\,
            I => \N__5704\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__5704\,
            I => \N__5701\
        );

    \I__1080\ : Odrv4
    port map (
            O => \N__5701\,
            I => \uart_tx_inst.n25\
        );

    \I__1079\ : InMux
    port map (
            O => \N__5698\,
            I => \uart_tx_inst.n1556\
        );

    \I__1078\ : InMux
    port map (
            O => \N__5695\,
            I => \N__5692\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__5692\,
            I => \N__5688\
        );

    \I__1076\ : InMux
    port map (
            O => \N__5691\,
            I => \N__5685\
        );

    \I__1075\ : Odrv4
    port map (
            O => \N__5688\,
            I => \uart_tx_inst.prescale_reg_12\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__5685\,
            I => \uart_tx_inst.prescale_reg_12\
        );

    \I__1073\ : InMux
    port map (
            O => \N__5680\,
            I => \N__5677\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__5677\,
            I => \N__5674\
        );

    \I__1071\ : Odrv4
    port map (
            O => \N__5674\,
            I => \uart_tx_inst.n24\
        );

    \I__1070\ : InMux
    port map (
            O => \N__5671\,
            I => \uart_tx_inst.n1557\
        );

    \I__1069\ : CascadeMux
    port map (
            O => \N__5668\,
            I => \N__5665\
        );

    \I__1068\ : InMux
    port map (
            O => \N__5665\,
            I => \N__5662\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__5662\,
            I => \N__5659\
        );

    \I__1066\ : Span4Mux_s2_h
    port map (
            O => \N__5659\,
            I => \N__5655\
        );

    \I__1065\ : InMux
    port map (
            O => \N__5658\,
            I => \N__5652\
        );

    \I__1064\ : Odrv4
    port map (
            O => \N__5655\,
            I => \uart_tx_inst.prescale_reg_13\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__5652\,
            I => \uart_tx_inst.prescale_reg_13\
        );

    \I__1062\ : InMux
    port map (
            O => \N__5647\,
            I => \N__5644\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__5644\,
            I => \N__5641\
        );

    \I__1060\ : Span4Mux_s2_v
    port map (
            O => \N__5641\,
            I => \N__5638\
        );

    \I__1059\ : Odrv4
    port map (
            O => \N__5638\,
            I => \uart_tx_inst.n23\
        );

    \I__1058\ : InMux
    port map (
            O => \N__5635\,
            I => \uart_tx_inst.n1558\
        );

    \I__1057\ : CascadeMux
    port map (
            O => \N__5632\,
            I => \uart_tx_inst.n860_cascade_\
        );

    \I__1056\ : InMux
    port map (
            O => \N__5629\,
            I => \bfn_11_2_0_\
        );

    \I__1055\ : InMux
    port map (
            O => \N__5626\,
            I => \N__5622\
        );

    \I__1054\ : InMux
    port map (
            O => \N__5625\,
            I => \N__5619\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__5622\,
            I => \uart_tx_inst.prescale_reg_1\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__5619\,
            I => \uart_tx_inst.prescale_reg_1\
        );

    \I__1051\ : InMux
    port map (
            O => \N__5614\,
            I => \uart_tx_inst.n1546\
        );

    \I__1050\ : InMux
    port map (
            O => \N__5611\,
            I => \N__5607\
        );

    \I__1049\ : InMux
    port map (
            O => \N__5610\,
            I => \N__5604\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__5607\,
            I => \uart_tx_inst.prescale_reg_2\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__5604\,
            I => \uart_tx_inst.prescale_reg_2\
        );

    \I__1046\ : InMux
    port map (
            O => \N__5599\,
            I => \uart_tx_inst.n1547\
        );

    \I__1045\ : SRMux
    port map (
            O => \N__5596\,
            I => \N__5593\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__5593\,
            I => \N__5590\
        );

    \I__1043\ : Odrv12
    port map (
            O => \N__5590\,
            I => \uart_tx_inst.n1170\
        );

    \I__1042\ : InMux
    port map (
            O => \N__5587\,
            I => \N__5583\
        );

    \I__1041\ : InMux
    port map (
            O => \N__5586\,
            I => \N__5580\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__5583\,
            I => \N__5577\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__5580\,
            I => \uart_tx_inst.prescale_reg_3\
        );

    \I__1038\ : Odrv4
    port map (
            O => \N__5577\,
            I => \uart_tx_inst.prescale_reg_3\
        );

    \I__1037\ : InMux
    port map (
            O => \N__5572\,
            I => \N__5569\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__5569\,
            I => \uart_tx_inst.n33\
        );

    \I__1035\ : InMux
    port map (
            O => \N__5566\,
            I => \uart_tx_inst.n1548\
        );

    \I__1034\ : InMux
    port map (
            O => \N__5563\,
            I => \uart_tx_inst.n1549\
        );

    \I__1033\ : InMux
    port map (
            O => \N__5560\,
            I => \uart_tx_inst.n1550\
        );

    \I__1032\ : InMux
    port map (
            O => \N__5557\,
            I => \N__5554\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__5554\,
            I => \N__5549\
        );

    \I__1030\ : InMux
    port map (
            O => \N__5553\,
            I => \N__5544\
        );

    \I__1029\ : InMux
    port map (
            O => \N__5552\,
            I => \N__5544\
        );

    \I__1028\ : Odrv4
    port map (
            O => \N__5549\,
            I => data_reg_4
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__5544\,
            I => data_reg_4
        );

    \I__1026\ : IoInMux
    port map (
            O => \N__5539\,
            I => \N__5536\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__5536\,
            I => \N__5533\
        );

    \I__1024\ : Span4Mux_s1_v
    port map (
            O => \N__5533\,
            I => \N__5530\
        );

    \I__1023\ : Odrv4
    port map (
            O => \N__5530\,
            I => output_axis_tdata_c_4
        );

    \I__1022\ : InMux
    port map (
            O => \N__5527\,
            I => \N__5523\
        );

    \I__1021\ : CascadeMux
    port map (
            O => \N__5526\,
            I => \N__5520\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__5523\,
            I => \N__5516\
        );

    \I__1019\ : InMux
    port map (
            O => \N__5520\,
            I => \N__5511\
        );

    \I__1018\ : InMux
    port map (
            O => \N__5519\,
            I => \N__5511\
        );

    \I__1017\ : Odrv12
    port map (
            O => \N__5516\,
            I => data_reg_5
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__5511\,
            I => data_reg_5
        );

    \I__1015\ : IoInMux
    port map (
            O => \N__5506\,
            I => \N__5503\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__5503\,
            I => \N__5500\
        );

    \I__1013\ : Span4Mux_s1_v
    port map (
            O => \N__5500\,
            I => \N__5497\
        );

    \I__1012\ : Odrv4
    port map (
            O => \N__5497\,
            I => output_axis_tdata_c_5
        );

    \I__1011\ : CascadeMux
    port map (
            O => \N__5494\,
            I => \N__5490\
        );

    \I__1010\ : InMux
    port map (
            O => \N__5493\,
            I => \N__5487\
        );

    \I__1009\ : InMux
    port map (
            O => \N__5490\,
            I => \N__5484\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__5487\,
            I => \N__5480\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__5484\,
            I => \N__5477\
        );

    \I__1006\ : InMux
    port map (
            O => \N__5483\,
            I => \N__5474\
        );

    \I__1005\ : Odrv12
    port map (
            O => \N__5480\,
            I => data_reg_1
        );

    \I__1004\ : Odrv4
    port map (
            O => \N__5477\,
            I => data_reg_1
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__5474\,
            I => data_reg_1
        );

    \I__1002\ : IoInMux
    port map (
            O => \N__5467\,
            I => \N__5464\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__5464\,
            I => \N__5461\
        );

    \I__1000\ : Span4Mux_s3_v
    port map (
            O => \N__5461\,
            I => \N__5458\
        );

    \I__999\ : Odrv4
    port map (
            O => \N__5458\,
            I => output_axis_tdata_c_1
        );

    \I__998\ : CascadeMux
    port map (
            O => \N__5455\,
            I => \N__5450\
        );

    \I__997\ : InMux
    port map (
            O => \N__5454\,
            I => \N__5447\
        );

    \I__996\ : InMux
    port map (
            O => \N__5453\,
            I => \N__5444\
        );

    \I__995\ : InMux
    port map (
            O => \N__5450\,
            I => \N__5441\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__5447\,
            I => \N__5438\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__5444\,
            I => data_reg_3
        );

    \I__992\ : LocalMux
    port map (
            O => \N__5441\,
            I => data_reg_3
        );

    \I__991\ : Odrv12
    port map (
            O => \N__5438\,
            I => data_reg_3
        );

    \I__990\ : IoInMux
    port map (
            O => \N__5431\,
            I => \N__5428\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__5428\,
            I => \N__5425\
        );

    \I__988\ : Span4Mux_s3_v
    port map (
            O => \N__5425\,
            I => \N__5422\
        );

    \I__987\ : Odrv4
    port map (
            O => \N__5422\,
            I => output_axis_tdata_c_3
        );

    \I__986\ : CEMux
    port map (
            O => \N__5419\,
            I => \N__5415\
        );

    \I__985\ : CEMux
    port map (
            O => \N__5418\,
            I => \N__5412\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__5415\,
            I => \N__5409\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__5412\,
            I => \N__5405\
        );

    \I__982\ : Span4Mux_v
    port map (
            O => \N__5409\,
            I => \N__5402\
        );

    \I__981\ : CEMux
    port map (
            O => \N__5408\,
            I => \N__5399\
        );

    \I__980\ : Span4Mux_v
    port map (
            O => \N__5405\,
            I => \N__5396\
        );

    \I__979\ : Span4Mux_s1_v
    port map (
            O => \N__5402\,
            I => \N__5393\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__5399\,
            I => \N__5390\
        );

    \I__977\ : Span4Mux_s1_v
    port map (
            O => \N__5396\,
            I => \N__5387\
        );

    \I__976\ : Odrv4
    port map (
            O => \N__5393\,
            I => n703
        );

    \I__975\ : Odrv12
    port map (
            O => \N__5390\,
            I => n703
        );

    \I__974\ : Odrv4
    port map (
            O => \N__5387\,
            I => n703
        );

    \I__973\ : CascadeMux
    port map (
            O => \N__5380\,
            I => \uart_tx_inst.n905_cascade_\
        );

    \I__972\ : CascadeMux
    port map (
            O => \N__5377\,
            I => \uart_tx_inst.n890_cascade_\
        );

    \I__971\ : InMux
    port map (
            O => \N__5374\,
            I => \N__5371\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__5371\,
            I => \N__5368\
        );

    \I__969\ : Odrv4
    port map (
            O => \N__5368\,
            I => \uart_tx_inst.n33_adj_198\
        );

    \I__968\ : InMux
    port map (
            O => \N__5365\,
            I => \N__5356\
        );

    \I__967\ : InMux
    port map (
            O => \N__5364\,
            I => \N__5348\
        );

    \I__966\ : InMux
    port map (
            O => \N__5363\,
            I => \N__5348\
        );

    \I__965\ : InMux
    port map (
            O => \N__5362\,
            I => \N__5348\
        );

    \I__964\ : InMux
    port map (
            O => \N__5361\,
            I => \N__5341\
        );

    \I__963\ : InMux
    port map (
            O => \N__5360\,
            I => \N__5341\
        );

    \I__962\ : InMux
    port map (
            O => \N__5359\,
            I => \N__5341\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__5356\,
            I => \N__5338\
        );

    \I__960\ : InMux
    port map (
            O => \N__5355\,
            I => \N__5335\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__5348\,
            I => n1711
        );

    \I__958\ : LocalMux
    port map (
            O => \N__5341\,
            I => n1711
        );

    \I__957\ : Odrv4
    port map (
            O => \N__5338\,
            I => n1711
        );

    \I__956\ : LocalMux
    port map (
            O => \N__5335\,
            I => n1711
        );

    \I__955\ : InMux
    port map (
            O => \N__5326\,
            I => \N__5317\
        );

    \I__954\ : InMux
    port map (
            O => \N__5325\,
            I => \N__5304\
        );

    \I__953\ : InMux
    port map (
            O => \N__5324\,
            I => \N__5304\
        );

    \I__952\ : InMux
    port map (
            O => \N__5323\,
            I => \N__5304\
        );

    \I__951\ : InMux
    port map (
            O => \N__5322\,
            I => \N__5304\
        );

    \I__950\ : InMux
    port map (
            O => \N__5321\,
            I => \N__5304\
        );

    \I__949\ : InMux
    port map (
            O => \N__5320\,
            I => \N__5304\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__5317\,
            I => \N__5301\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__5304\,
            I => n1220
        );

    \I__946\ : Odrv4
    port map (
            O => \N__5301\,
            I => n1220
        );

    \I__945\ : InMux
    port map (
            O => \N__5296\,
            I => \N__5286\
        );

    \I__944\ : InMux
    port map (
            O => \N__5295\,
            I => \N__5286\
        );

    \I__943\ : InMux
    port map (
            O => \N__5294\,
            I => \N__5283\
        );

    \I__942\ : InMux
    port map (
            O => \N__5293\,
            I => \N__5279\
        );

    \I__941\ : InMux
    port map (
            O => \N__5292\,
            I => \N__5276\
        );

    \I__940\ : InMux
    port map (
            O => \N__5291\,
            I => \N__5273\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__5286\,
            I => \N__5266\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__5283\,
            I => \N__5263\
        );

    \I__937\ : InMux
    port map (
            O => \N__5282\,
            I => \N__5260\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__5279\,
            I => \N__5257\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__5276\,
            I => \N__5254\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__5273\,
            I => \N__5251\
        );

    \I__933\ : InMux
    port map (
            O => \N__5272\,
            I => \N__5242\
        );

    \I__932\ : InMux
    port map (
            O => \N__5271\,
            I => \N__5242\
        );

    \I__931\ : InMux
    port map (
            O => \N__5270\,
            I => \N__5242\
        );

    \I__930\ : InMux
    port map (
            O => \N__5269\,
            I => \N__5242\
        );

    \I__929\ : Span4Mux_v
    port map (
            O => \N__5266\,
            I => \N__5233\
        );

    \I__928\ : Span4Mux_h
    port map (
            O => \N__5263\,
            I => \N__5233\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__5260\,
            I => \N__5233\
        );

    \I__926\ : Span4Mux_v
    port map (
            O => \N__5257\,
            I => \N__5233\
        );

    \I__925\ : Span12Mux_v
    port map (
            O => \N__5254\,
            I => \N__5230\
        );

    \I__924\ : Span12Mux_s7_h
    port map (
            O => \N__5251\,
            I => \N__5225\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__5242\,
            I => \N__5225\
        );

    \I__922\ : Odrv4
    port map (
            O => \N__5233\,
            I => rxd_reg
        );

    \I__921\ : Odrv12
    port map (
            O => \N__5230\,
            I => rxd_reg
        );

    \I__920\ : Odrv12
    port map (
            O => \N__5225\,
            I => rxd_reg
        );

    \I__919\ : IoInMux
    port map (
            O => \N__5218\,
            I => \N__5215\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__5215\,
            I => \N__5212\
        );

    \I__917\ : Span4Mux_s3_h
    port map (
            O => \N__5212\,
            I => \N__5209\
        );

    \I__916\ : Odrv4
    port map (
            O => \N__5209\,
            I => rx_frame_error_c
        );

    \I__915\ : SRMux
    port map (
            O => \N__5206\,
            I => \N__5203\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__5203\,
            I => \N__5200\
        );

    \I__913\ : Span4Mux_h
    port map (
            O => \N__5200\,
            I => \N__5197\
        );

    \I__912\ : Odrv4
    port map (
            O => \N__5197\,
            I => n697
        );

    \I__911\ : InMux
    port map (
            O => \N__5194\,
            I => \N__5190\
        );

    \I__910\ : CascadeMux
    port map (
            O => \N__5193\,
            I => \N__5187\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__5190\,
            I => \N__5183\
        );

    \I__908\ : InMux
    port map (
            O => \N__5187\,
            I => \N__5178\
        );

    \I__907\ : InMux
    port map (
            O => \N__5186\,
            I => \N__5178\
        );

    \I__906\ : Odrv4
    port map (
            O => \N__5183\,
            I => data_reg_6
        );

    \I__905\ : LocalMux
    port map (
            O => \N__5178\,
            I => data_reg_6
        );

    \I__904\ : IoInMux
    port map (
            O => \N__5173\,
            I => \N__5170\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__5170\,
            I => \N__5167\
        );

    \I__902\ : Odrv12
    port map (
            O => \N__5167\,
            I => output_axis_tdata_c_6
        );

    \I__901\ : CascadeMux
    port map (
            O => \N__5164\,
            I => \N__5159\
        );

    \I__900\ : CascadeMux
    port map (
            O => \N__5163\,
            I => \N__5156\
        );

    \I__899\ : InMux
    port map (
            O => \N__5162\,
            I => \N__5153\
        );

    \I__898\ : InMux
    port map (
            O => \N__5159\,
            I => \N__5150\
        );

    \I__897\ : InMux
    port map (
            O => \N__5156\,
            I => \N__5147\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__5153\,
            I => \N__5144\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__5150\,
            I => data_reg_2
        );

    \I__894\ : LocalMux
    port map (
            O => \N__5147\,
            I => data_reg_2
        );

    \I__893\ : Odrv12
    port map (
            O => \N__5144\,
            I => data_reg_2
        );

    \I__892\ : IoInMux
    port map (
            O => \N__5137\,
            I => \N__5134\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__5134\,
            I => \N__5131\
        );

    \I__890\ : IoSpan4Mux
    port map (
            O => \N__5131\,
            I => \N__5128\
        );

    \I__889\ : Span4Mux_s1_v
    port map (
            O => \N__5128\,
            I => \N__5125\
        );

    \I__888\ : Odrv4
    port map (
            O => \N__5125\,
            I => output_axis_tdata_c_2
        );

    \I__887\ : InMux
    port map (
            O => \N__5122\,
            I => \N__5119\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__5119\,
            I => \N__5115\
        );

    \I__885\ : CascadeMux
    port map (
            O => \N__5118\,
            I => \N__5112\
        );

    \I__884\ : Span4Mux_v
    port map (
            O => \N__5115\,
            I => \N__5108\
        );

    \I__883\ : InMux
    port map (
            O => \N__5112\,
            I => \N__5105\
        );

    \I__882\ : InMux
    port map (
            O => \N__5111\,
            I => \N__5102\
        );

    \I__881\ : Odrv4
    port map (
            O => \N__5108\,
            I => data_reg_7
        );

    \I__880\ : LocalMux
    port map (
            O => \N__5105\,
            I => data_reg_7
        );

    \I__879\ : LocalMux
    port map (
            O => \N__5102\,
            I => data_reg_7
        );

    \I__878\ : IoInMux
    port map (
            O => \N__5095\,
            I => \N__5092\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__5092\,
            I => \N__5089\
        );

    \I__876\ : Odrv12
    port map (
            O => \N__5089\,
            I => output_axis_tdata_c_7
        );

    \I__875\ : InMux
    port map (
            O => \N__5086\,
            I => \N__5083\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__5083\,
            I => \N__5080\
        );

    \I__873\ : Odrv4
    port map (
            O => \N__5080\,
            I => \uart_rx_inst.n1750\
        );

    \I__872\ : InMux
    port map (
            O => \N__5077\,
            I => \N__5074\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__5074\,
            I => \N__5071\
        );

    \I__870\ : Odrv4
    port map (
            O => \N__5071\,
            I => \uart_rx_inst.n1755\
        );

    \I__869\ : CascadeMux
    port map (
            O => \N__5068\,
            I => \N__5065\
        );

    \I__868\ : InMux
    port map (
            O => \N__5065\,
            I => \N__5062\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__5062\,
            I => \uart_rx_inst.n1754\
        );

    \I__866\ : InMux
    port map (
            O => \N__5059\,
            I => \N__5056\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__5056\,
            I => \N__5053\
        );

    \I__864\ : Odrv4
    port map (
            O => \N__5053\,
            I => \uart_rx_inst.n1751\
        );

    \I__863\ : InMux
    port map (
            O => \N__5050\,
            I => \N__5047\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__5047\,
            I => \N__5044\
        );

    \I__861\ : Odrv4
    port map (
            O => \N__5044\,
            I => \uart_rx_inst.n1758\
        );

    \I__860\ : InMux
    port map (
            O => \N__5041\,
            I => \N__5038\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__5038\,
            I => \uart_rx_inst.n1742\
        );

    \I__858\ : InMux
    port map (
            O => \N__5035\,
            I => \N__5032\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__5032\,
            I => \N__5029\
        );

    \I__856\ : Odrv12
    port map (
            O => \N__5029\,
            I => \uart_rx_inst.n1739\
        );

    \I__855\ : InMux
    port map (
            O => \N__5026\,
            I => \N__5023\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__5023\,
            I => \N__5020\
        );

    \I__853\ : Odrv12
    port map (
            O => \N__5020\,
            I => \uart_rx_inst.n1757\
        );

    \I__852\ : CascadeMux
    port map (
            O => \N__5017\,
            I => \N__5014\
        );

    \I__851\ : InMux
    port map (
            O => \N__5014\,
            I => \N__5010\
        );

    \I__850\ : InMux
    port map (
            O => \N__5013\,
            I => \N__5007\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__5010\,
            I => \uart_rx_inst.prescale_reg_15\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__5007\,
            I => \uart_rx_inst.prescale_reg_15\
        );

    \I__847\ : InMux
    port map (
            O => \N__5002\,
            I => \N__4999\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__4999\,
            I => \uart_rx_inst.n749\
        );

    \I__845\ : InMux
    port map (
            O => \N__4996\,
            I => \uart_rx_inst.n1578\
        );

    \I__844\ : CascadeMux
    port map (
            O => \N__4993\,
            I => \N__4989\
        );

    \I__843\ : InMux
    port map (
            O => \N__4992\,
            I => \N__4986\
        );

    \I__842\ : InMux
    port map (
            O => \N__4989\,
            I => \N__4983\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__4986\,
            I => \uart_rx_inst.prescale_reg_16\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__4983\,
            I => \uart_rx_inst.prescale_reg_16\
        );

    \I__839\ : InMux
    port map (
            O => \N__4978\,
            I => \N__4975\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__4975\,
            I => \uart_rx_inst.n744\
        );

    \I__837\ : InMux
    port map (
            O => \N__4972\,
            I => \bfn_9_7_0_\
        );

    \I__836\ : CascadeMux
    port map (
            O => \N__4969\,
            I => \N__4966\
        );

    \I__835\ : InMux
    port map (
            O => \N__4966\,
            I => \N__4963\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__4963\,
            I => \N__4959\
        );

    \I__833\ : InMux
    port map (
            O => \N__4962\,
            I => \N__4956\
        );

    \I__832\ : Odrv4
    port map (
            O => \N__4959\,
            I => \uart_rx_inst.prescale_reg_17\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__4956\,
            I => \uart_rx_inst.prescale_reg_17\
        );

    \I__830\ : InMux
    port map (
            O => \N__4951\,
            I => \N__4948\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__4948\,
            I => \uart_rx_inst.n739\
        );

    \I__828\ : InMux
    port map (
            O => \N__4945\,
            I => \uart_rx_inst.n1580\
        );

    \I__827\ : CascadeMux
    port map (
            O => \N__4942\,
            I => \N__4929\
        );

    \I__826\ : CascadeMux
    port map (
            O => \N__4941\,
            I => \N__4925\
        );

    \I__825\ : CascadeMux
    port map (
            O => \N__4940\,
            I => \N__4921\
        );

    \I__824\ : CascadeMux
    port map (
            O => \N__4939\,
            I => \N__4917\
        );

    \I__823\ : CascadeMux
    port map (
            O => \N__4938\,
            I => \N__4913\
        );

    \I__822\ : CascadeMux
    port map (
            O => \N__4937\,
            I => \N__4910\
        );

    \I__821\ : CascadeMux
    port map (
            O => \N__4936\,
            I => \N__4906\
        );

    \I__820\ : CascadeMux
    port map (
            O => \N__4935\,
            I => \N__4902\
        );

    \I__819\ : CascadeMux
    port map (
            O => \N__4934\,
            I => \N__4898\
        );

    \I__818\ : InMux
    port map (
            O => \N__4933\,
            I => \N__4891\
        );

    \I__817\ : InMux
    port map (
            O => \N__4932\,
            I => \N__4891\
        );

    \I__816\ : InMux
    port map (
            O => \N__4929\,
            I => \N__4891\
        );

    \I__815\ : InMux
    port map (
            O => \N__4928\,
            I => \N__4874\
        );

    \I__814\ : InMux
    port map (
            O => \N__4925\,
            I => \N__4874\
        );

    \I__813\ : InMux
    port map (
            O => \N__4924\,
            I => \N__4874\
        );

    \I__812\ : InMux
    port map (
            O => \N__4921\,
            I => \N__4874\
        );

    \I__811\ : InMux
    port map (
            O => \N__4920\,
            I => \N__4874\
        );

    \I__810\ : InMux
    port map (
            O => \N__4917\,
            I => \N__4874\
        );

    \I__809\ : InMux
    port map (
            O => \N__4916\,
            I => \N__4874\
        );

    \I__808\ : InMux
    port map (
            O => \N__4913\,
            I => \N__4874\
        );

    \I__807\ : InMux
    port map (
            O => \N__4910\,
            I => \N__4859\
        );

    \I__806\ : InMux
    port map (
            O => \N__4909\,
            I => \N__4859\
        );

    \I__805\ : InMux
    port map (
            O => \N__4906\,
            I => \N__4859\
        );

    \I__804\ : InMux
    port map (
            O => \N__4905\,
            I => \N__4859\
        );

    \I__803\ : InMux
    port map (
            O => \N__4902\,
            I => \N__4859\
        );

    \I__802\ : InMux
    port map (
            O => \N__4901\,
            I => \N__4859\
        );

    \I__801\ : InMux
    port map (
            O => \N__4898\,
            I => \N__4859\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__4891\,
            I => \uart_rx_inst.n712\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__4874\,
            I => \uart_rx_inst.n712\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__4859\,
            I => \uart_rx_inst.n712\
        );

    \I__797\ : InMux
    port map (
            O => \N__4852\,
            I => \N__4849\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__4849\,
            I => \N__4845\
        );

    \I__795\ : InMux
    port map (
            O => \N__4848\,
            I => \N__4842\
        );

    \I__794\ : Odrv4
    port map (
            O => \N__4845\,
            I => \uart_rx_inst.prescale_reg_18\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__4842\,
            I => \uart_rx_inst.prescale_reg_18\
        );

    \I__792\ : InMux
    port map (
            O => \N__4837\,
            I => \uart_rx_inst.n1581\
        );

    \I__791\ : InMux
    port map (
            O => \N__4834\,
            I => \N__4831\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__4831\,
            I => \N__4828\
        );

    \I__789\ : Odrv4
    port map (
            O => \N__4828\,
            I => \uart_rx_inst.n729\
        );

    \I__788\ : InMux
    port map (
            O => \N__4825\,
            I => \N__4822\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__4822\,
            I => \uart_rx_inst.n1743\
        );

    \I__786\ : InMux
    port map (
            O => \N__4819\,
            I => \N__4816\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__4816\,
            I => \uart_rx_inst.n1740\
        );

    \I__784\ : InMux
    port map (
            O => \N__4813\,
            I => \N__4810\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__4810\,
            I => \uart_rx_inst.n1741\
        );

    \I__782\ : InMux
    port map (
            O => \N__4807\,
            I => \N__4804\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__4804\,
            I => \uart_rx_inst.n1747\
        );

    \I__780\ : InMux
    port map (
            O => \N__4801\,
            I => \N__4798\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__4798\,
            I => \uart_rx_inst.n1745\
        );

    \I__778\ : InMux
    port map (
            O => \N__4795\,
            I => \N__4792\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__4792\,
            I => \N__4788\
        );

    \I__776\ : CascadeMux
    port map (
            O => \N__4791\,
            I => \N__4785\
        );

    \I__775\ : Span4Mux_v
    port map (
            O => \N__4788\,
            I => \N__4782\
        );

    \I__774\ : InMux
    port map (
            O => \N__4785\,
            I => \N__4779\
        );

    \I__773\ : Odrv4
    port map (
            O => \N__4782\,
            I => \uart_rx_inst.prescale_reg_8\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__4779\,
            I => \uart_rx_inst.prescale_reg_8\
        );

    \I__771\ : InMux
    port map (
            O => \N__4774\,
            I => \N__4771\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__4771\,
            I => \N__4768\
        );

    \I__769\ : Span4Mux_v
    port map (
            O => \N__4768\,
            I => \N__4765\
        );

    \I__768\ : Odrv4
    port map (
            O => \N__4765\,
            I => \uart_rx_inst.n784\
        );

    \I__767\ : InMux
    port map (
            O => \N__4762\,
            I => \bfn_9_6_0_\
        );

    \I__766\ : CascadeMux
    port map (
            O => \N__4759\,
            I => \N__4755\
        );

    \I__765\ : CascadeMux
    port map (
            O => \N__4758\,
            I => \N__4752\
        );

    \I__764\ : InMux
    port map (
            O => \N__4755\,
            I => \N__4749\
        );

    \I__763\ : InMux
    port map (
            O => \N__4752\,
            I => \N__4746\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__4749\,
            I => \N__4743\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__4746\,
            I => \uart_rx_inst.prescale_reg_9\
        );

    \I__760\ : Odrv4
    port map (
            O => \N__4743\,
            I => \uart_rx_inst.prescale_reg_9\
        );

    \I__759\ : InMux
    port map (
            O => \N__4738\,
            I => \N__4735\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__4735\,
            I => \uart_rx_inst.n779\
        );

    \I__757\ : InMux
    port map (
            O => \N__4732\,
            I => \uart_rx_inst.n1572\
        );

    \I__756\ : InMux
    port map (
            O => \N__4729\,
            I => \N__4726\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__4726\,
            I => \N__4723\
        );

    \I__754\ : Span4Mux_h
    port map (
            O => \N__4723\,
            I => \N__4720\
        );

    \I__753\ : Odrv4
    port map (
            O => \N__4720\,
            I => \uart_rx_inst.n1744\
        );

    \I__752\ : CascadeMux
    port map (
            O => \N__4717\,
            I => \N__4713\
        );

    \I__751\ : InMux
    port map (
            O => \N__4716\,
            I => \N__4710\
        );

    \I__750\ : InMux
    port map (
            O => \N__4713\,
            I => \N__4707\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__4710\,
            I => \uart_rx_inst.prescale_reg_10\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__4707\,
            I => \uart_rx_inst.prescale_reg_10\
        );

    \I__747\ : InMux
    port map (
            O => \N__4702\,
            I => \N__4699\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__4699\,
            I => \uart_rx_inst.n774\
        );

    \I__745\ : InMux
    port map (
            O => \N__4696\,
            I => \uart_rx_inst.n1573\
        );

    \I__744\ : CascadeMux
    port map (
            O => \N__4693\,
            I => \N__4690\
        );

    \I__743\ : InMux
    port map (
            O => \N__4690\,
            I => \N__4686\
        );

    \I__742\ : InMux
    port map (
            O => \N__4689\,
            I => \N__4683\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__4686\,
            I => \uart_rx_inst.prescale_reg_11\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__4683\,
            I => \uart_rx_inst.prescale_reg_11\
        );

    \I__739\ : InMux
    port map (
            O => \N__4678\,
            I => \N__4675\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__4675\,
            I => \uart_rx_inst.n769\
        );

    \I__737\ : InMux
    port map (
            O => \N__4672\,
            I => \uart_rx_inst.n1574\
        );

    \I__736\ : InMux
    port map (
            O => \N__4669\,
            I => \N__4665\
        );

    \I__735\ : InMux
    port map (
            O => \N__4668\,
            I => \N__4662\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__4665\,
            I => \uart_rx_inst.prescale_reg_12\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__4662\,
            I => \uart_rx_inst.prescale_reg_12\
        );

    \I__732\ : CascadeMux
    port map (
            O => \N__4657\,
            I => \N__4654\
        );

    \I__731\ : InMux
    port map (
            O => \N__4654\,
            I => \N__4651\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__4651\,
            I => \uart_rx_inst.n764\
        );

    \I__729\ : InMux
    port map (
            O => \N__4648\,
            I => \uart_rx_inst.n1575\
        );

    \I__728\ : CascadeMux
    port map (
            O => \N__4645\,
            I => \N__4642\
        );

    \I__727\ : InMux
    port map (
            O => \N__4642\,
            I => \N__4638\
        );

    \I__726\ : InMux
    port map (
            O => \N__4641\,
            I => \N__4635\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__4638\,
            I => \uart_rx_inst.prescale_reg_13\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__4635\,
            I => \uart_rx_inst.prescale_reg_13\
        );

    \I__723\ : InMux
    port map (
            O => \N__4630\,
            I => \N__4627\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__4627\,
            I => \uart_rx_inst.n759\
        );

    \I__721\ : InMux
    port map (
            O => \N__4624\,
            I => \uart_rx_inst.n1576\
        );

    \I__720\ : InMux
    port map (
            O => \N__4621\,
            I => \N__4618\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__4618\,
            I => \N__4614\
        );

    \I__718\ : InMux
    port map (
            O => \N__4617\,
            I => \N__4611\
        );

    \I__717\ : Odrv4
    port map (
            O => \N__4614\,
            I => \uart_rx_inst.prescale_reg_14\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__4611\,
            I => \uart_rx_inst.prescale_reg_14\
        );

    \I__715\ : InMux
    port map (
            O => \N__4606\,
            I => \N__4603\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__4603\,
            I => \uart_rx_inst.n754\
        );

    \I__713\ : InMux
    port map (
            O => \N__4600\,
            I => \uart_rx_inst.n1577\
        );

    \I__712\ : InMux
    port map (
            O => \N__4597\,
            I => \N__4591\
        );

    \I__711\ : InMux
    port map (
            O => \N__4596\,
            I => \N__4586\
        );

    \I__710\ : InMux
    port map (
            O => \N__4595\,
            I => \N__4586\
        );

    \I__709\ : InMux
    port map (
            O => \N__4594\,
            I => \N__4583\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__4591\,
            I => \uart_rx_inst.n509\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__4586\,
            I => \uart_rx_inst.n509\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__4583\,
            I => \uart_rx_inst.n509\
        );

    \I__705\ : CascadeMux
    port map (
            O => \N__4576\,
            I => \N__4572\
        );

    \I__704\ : InMux
    port map (
            O => \N__4575\,
            I => \N__4569\
        );

    \I__703\ : InMux
    port map (
            O => \N__4572\,
            I => \N__4566\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__4569\,
            I => \N__4563\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__4566\,
            I => \uart_rx_inst.prescale_reg_0\
        );

    \I__700\ : Odrv4
    port map (
            O => \N__4563\,
            I => \uart_rx_inst.prescale_reg_0\
        );

    \I__699\ : InMux
    port map (
            O => \N__4558\,
            I => \bfn_9_5_0_\
        );

    \I__698\ : CEMux
    port map (
            O => \N__4555\,
            I => \N__4552\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__4552\,
            I => \N__4549\
        );

    \I__696\ : Span4Mux_v
    port map (
            O => \N__4549\,
            I => \N__4546\
        );

    \I__695\ : Odrv4
    port map (
            O => \N__4546\,
            I => \uart_rx_inst.n1648\
        );

    \I__694\ : SRMux
    port map (
            O => \N__4543\,
            I => \N__4540\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__4540\,
            I => \N__4537\
        );

    \I__692\ : Span4Mux_s3_h
    port map (
            O => \N__4537\,
            I => \N__4534\
        );

    \I__691\ : Span4Mux_v
    port map (
            O => \N__4534\,
            I => \N__4531\
        );

    \I__690\ : Odrv4
    port map (
            O => \N__4531\,
            I => \uart_rx_inst.n1141\
        );

    \I__689\ : InMux
    port map (
            O => \N__4528\,
            I => \N__4525\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__4525\,
            I => \N__4522\
        );

    \I__687\ : Span4Mux_s3_h
    port map (
            O => \N__4522\,
            I => \N__4518\
        );

    \I__686\ : InMux
    port map (
            O => \N__4521\,
            I => \N__4515\
        );

    \I__685\ : Odrv4
    port map (
            O => \N__4518\,
            I => \uart_rx_inst.prescale_reg_1\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__4515\,
            I => \uart_rx_inst.prescale_reg_1\
        );

    \I__683\ : InMux
    port map (
            O => \N__4510\,
            I => \N__4507\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__4507\,
            I => \N__4504\
        );

    \I__681\ : Odrv4
    port map (
            O => \N__4504\,
            I => \uart_rx_inst.n819\
        );

    \I__680\ : InMux
    port map (
            O => \N__4501\,
            I => \uart_rx_inst.n1564\
        );

    \I__679\ : CascadeMux
    port map (
            O => \N__4498\,
            I => \N__4495\
        );

    \I__678\ : InMux
    port map (
            O => \N__4495\,
            I => \N__4492\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__4492\,
            I => \N__4489\
        );

    \I__676\ : Span4Mux_h
    port map (
            O => \N__4489\,
            I => \N__4485\
        );

    \I__675\ : InMux
    port map (
            O => \N__4488\,
            I => \N__4482\
        );

    \I__674\ : Odrv4
    port map (
            O => \N__4485\,
            I => \uart_rx_inst.prescale_reg_2\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__4482\,
            I => \uart_rx_inst.prescale_reg_2\
        );

    \I__672\ : InMux
    port map (
            O => \N__4477\,
            I => \N__4474\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__4474\,
            I => \N__4471\
        );

    \I__670\ : Span4Mux_v
    port map (
            O => \N__4471\,
            I => \N__4468\
        );

    \I__669\ : Odrv4
    port map (
            O => \N__4468\,
            I => \uart_rx_inst.n814\
        );

    \I__668\ : InMux
    port map (
            O => \N__4465\,
            I => \uart_rx_inst.n1565\
        );

    \I__667\ : InMux
    port map (
            O => \N__4462\,
            I => \N__4458\
        );

    \I__666\ : InMux
    port map (
            O => \N__4461\,
            I => \N__4455\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__4458\,
            I => \uart_rx_inst.prescale_reg_3\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__4455\,
            I => \uart_rx_inst.prescale_reg_3\
        );

    \I__663\ : InMux
    port map (
            O => \N__4450\,
            I => \N__4447\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__4447\,
            I => \uart_rx_inst.n809\
        );

    \I__661\ : InMux
    port map (
            O => \N__4444\,
            I => \uart_rx_inst.n1566\
        );

    \I__660\ : CascadeMux
    port map (
            O => \N__4441\,
            I => \N__4438\
        );

    \I__659\ : InMux
    port map (
            O => \N__4438\,
            I => \N__4435\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__4435\,
            I => \N__4431\
        );

    \I__657\ : InMux
    port map (
            O => \N__4434\,
            I => \N__4428\
        );

    \I__656\ : Odrv4
    port map (
            O => \N__4431\,
            I => \uart_rx_inst.prescale_reg_4\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__4428\,
            I => \uart_rx_inst.prescale_reg_4\
        );

    \I__654\ : InMux
    port map (
            O => \N__4423\,
            I => \N__4420\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__4420\,
            I => \N__4417\
        );

    \I__652\ : Odrv4
    port map (
            O => \N__4417\,
            I => \uart_rx_inst.n804\
        );

    \I__651\ : InMux
    port map (
            O => \N__4414\,
            I => \uart_rx_inst.n1567\
        );

    \I__650\ : InMux
    port map (
            O => \N__4411\,
            I => \N__4408\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__4408\,
            I => \N__4405\
        );

    \I__648\ : Span4Mux_h
    port map (
            O => \N__4405\,
            I => \N__4402\
        );

    \I__647\ : Odrv4
    port map (
            O => \N__4402\,
            I => \uart_rx_inst.n1756\
        );

    \I__646\ : InMux
    port map (
            O => \N__4399\,
            I => \N__4396\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__4396\,
            I => \N__4392\
        );

    \I__644\ : InMux
    port map (
            O => \N__4395\,
            I => \N__4389\
        );

    \I__643\ : Odrv4
    port map (
            O => \N__4392\,
            I => \uart_rx_inst.prescale_reg_5\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__4389\,
            I => \uart_rx_inst.prescale_reg_5\
        );

    \I__641\ : InMux
    port map (
            O => \N__4384\,
            I => \N__4381\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__4381\,
            I => \N__4378\
        );

    \I__639\ : Odrv4
    port map (
            O => \N__4378\,
            I => \uart_rx_inst.n799\
        );

    \I__638\ : InMux
    port map (
            O => \N__4375\,
            I => \uart_rx_inst.n1568\
        );

    \I__637\ : CascadeMux
    port map (
            O => \N__4372\,
            I => \N__4369\
        );

    \I__636\ : InMux
    port map (
            O => \N__4369\,
            I => \N__4365\
        );

    \I__635\ : InMux
    port map (
            O => \N__4368\,
            I => \N__4362\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__4365\,
            I => \uart_rx_inst.prescale_reg_6\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__4362\,
            I => \uart_rx_inst.prescale_reg_6\
        );

    \I__632\ : InMux
    port map (
            O => \N__4357\,
            I => \N__4354\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__4354\,
            I => \uart_rx_inst.n794\
        );

    \I__630\ : InMux
    port map (
            O => \N__4351\,
            I => \uart_rx_inst.n1569\
        );

    \I__629\ : InMux
    port map (
            O => \N__4348\,
            I => \N__4344\
        );

    \I__628\ : InMux
    port map (
            O => \N__4347\,
            I => \N__4341\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__4344\,
            I => \uart_rx_inst.prescale_reg_7\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__4341\,
            I => \uart_rx_inst.prescale_reg_7\
        );

    \I__625\ : InMux
    port map (
            O => \N__4336\,
            I => \N__4333\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__4333\,
            I => \uart_rx_inst.n789\
        );

    \I__623\ : InMux
    port map (
            O => \N__4330\,
            I => \uart_rx_inst.n1570\
        );

    \I__622\ : CascadeMux
    port map (
            O => \N__4327\,
            I => \uart_tx_inst.n880_cascade_\
        );

    \I__621\ : CascadeMux
    port map (
            O => \N__4324\,
            I => \uart_tx_inst.n895_cascade_\
        );

    \I__620\ : CascadeMux
    port map (
            O => \N__4321\,
            I => \uart_tx_inst.n900_cascade_\
        );

    \I__619\ : InMux
    port map (
            O => \N__4318\,
            I => \N__4315\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__4315\,
            I => \uart_tx_inst.n925\
        );

    \I__617\ : InMux
    port map (
            O => \N__4312\,
            I => \N__4309\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__4309\,
            I => \uart_tx_inst.n935\
        );

    \I__615\ : CascadeMux
    port map (
            O => \N__4306\,
            I => \uart_tx_inst.n920_cascade_\
        );

    \I__614\ : CascadeMux
    port map (
            O => \N__4303\,
            I => \uart_tx_inst.n930_cascade_\
        );

    \I__613\ : InMux
    port map (
            O => \N__4300\,
            I => \N__4297\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__4297\,
            I => \uart_tx_inst.n31_adj_199\
        );

    \I__611\ : InMux
    port map (
            O => \N__4294\,
            I => \N__4291\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__4291\,
            I => \uart_tx_inst.n915\
        );

    \I__609\ : CascadeMux
    port map (
            O => \N__4288\,
            I => \uart_tx_inst.n875_cascade_\
        );

    \I__608\ : SRMux
    port map (
            O => \N__4285\,
            I => \N__4282\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__4282\,
            I => \N__4279\
        );

    \I__606\ : Span4Mux_h
    port map (
            O => \N__4279\,
            I => \N__4276\
        );

    \I__605\ : Odrv4
    port map (
            O => \N__4276\,
            I => n1167
        );

    \I__604\ : InMux
    port map (
            O => \N__4273\,
            I => \N__4265\
        );

    \I__603\ : InMux
    port map (
            O => \N__4272\,
            I => \N__4265\
        );

    \I__602\ : InMux
    port map (
            O => \N__4271\,
            I => \N__4258\
        );

    \I__601\ : CascadeMux
    port map (
            O => \N__4270\,
            I => \N__4254\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__4265\,
            I => \N__4250\
        );

    \I__599\ : InMux
    port map (
            O => \N__4264\,
            I => \N__4247\
        );

    \I__598\ : InMux
    port map (
            O => \N__4263\,
            I => \N__4242\
        );

    \I__597\ : InMux
    port map (
            O => \N__4262\,
            I => \N__4242\
        );

    \I__596\ : InMux
    port map (
            O => \N__4261\,
            I => \N__4239\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__4258\,
            I => \N__4236\
        );

    \I__594\ : InMux
    port map (
            O => \N__4257\,
            I => \N__4229\
        );

    \I__593\ : InMux
    port map (
            O => \N__4254\,
            I => \N__4229\
        );

    \I__592\ : InMux
    port map (
            O => \N__4253\,
            I => \N__4229\
        );

    \I__591\ : Span4Mux_v
    port map (
            O => \N__4250\,
            I => \N__4226\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__4247\,
            I => bit_cnt_0
        );

    \I__589\ : LocalMux
    port map (
            O => \N__4242\,
            I => bit_cnt_0
        );

    \I__588\ : LocalMux
    port map (
            O => \N__4239\,
            I => bit_cnt_0
        );

    \I__587\ : Odrv4
    port map (
            O => \N__4236\,
            I => bit_cnt_0
        );

    \I__586\ : LocalMux
    port map (
            O => \N__4229\,
            I => bit_cnt_0
        );

    \I__585\ : Odrv4
    port map (
            O => \N__4226\,
            I => bit_cnt_0
        );

    \I__584\ : InMux
    port map (
            O => \N__4213\,
            I => \N__4207\
        );

    \I__583\ : InMux
    port map (
            O => \N__4212\,
            I => \N__4201\
        );

    \I__582\ : InMux
    port map (
            O => \N__4211\,
            I => \N__4201\
        );

    \I__581\ : InMux
    port map (
            O => \N__4210\,
            I => \N__4198\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__4207\,
            I => \N__4195\
        );

    \I__579\ : InMux
    port map (
            O => \N__4206\,
            I => \N__4192\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__4201\,
            I => \N__4189\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__4198\,
            I => \uart_rx_inst.n677\
        );

    \I__576\ : Odrv4
    port map (
            O => \N__4195\,
            I => \uart_rx_inst.n677\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__4192\,
            I => \uart_rx_inst.n677\
        );

    \I__574\ : Odrv4
    port map (
            O => \N__4189\,
            I => \uart_rx_inst.n677\
        );

    \I__573\ : CascadeMux
    port map (
            O => \N__4180\,
            I => \N__4177\
        );

    \I__572\ : InMux
    port map (
            O => \N__4177\,
            I => \N__4174\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__4174\,
            I => \N__4170\
        );

    \I__570\ : InMux
    port map (
            O => \N__4173\,
            I => \N__4167\
        );

    \I__569\ : Odrv4
    port map (
            O => \N__4170\,
            I => \uart_rx_inst.output_axis_tvalid_N_172\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__4167\,
            I => \uart_rx_inst.output_axis_tvalid_N_172\
        );

    \I__567\ : InMux
    port map (
            O => \N__4162\,
            I => \N__4156\
        );

    \I__566\ : InMux
    port map (
            O => \N__4161\,
            I => \N__4149\
        );

    \I__565\ : InMux
    port map (
            O => \N__4160\,
            I => \N__4149\
        );

    \I__564\ : InMux
    port map (
            O => \N__4159\,
            I => \N__4149\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__4156\,
            I => \uart_rx_inst.output_axis_tvalid_N_173\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__4149\,
            I => \uart_rx_inst.output_axis_tvalid_N_173\
        );

    \I__561\ : CascadeMux
    port map (
            O => \N__4144\,
            I => \n695_cascade_\
        );

    \I__560\ : InMux
    port map (
            O => \N__4141\,
            I => \N__4138\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__4138\,
            I => n695
        );

    \I__558\ : InMux
    port map (
            O => \N__4135\,
            I => \N__4131\
        );

    \I__557\ : InMux
    port map (
            O => \N__4134\,
            I => \N__4128\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__4131\,
            I => \N__4120\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__4128\,
            I => \N__4120\
        );

    \I__554\ : InMux
    port map (
            O => \N__4127\,
            I => \N__4117\
        );

    \I__553\ : InMux
    port map (
            O => \N__4126\,
            I => \N__4114\
        );

    \I__552\ : InMux
    port map (
            O => \N__4125\,
            I => \N__4111\
        );

    \I__551\ : Span4Mux_v
    port map (
            O => \N__4120\,
            I => \N__4104\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__4117\,
            I => \N__4104\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__4114\,
            I => \N__4104\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__4111\,
            I => \output_axis_tvalid_N_175\
        );

    \I__547\ : Odrv4
    port map (
            O => \N__4104\,
            I => \output_axis_tvalid_N_175\
        );

    \I__546\ : InMux
    port map (
            O => \N__4099\,
            I => \N__4095\
        );

    \I__545\ : InMux
    port map (
            O => \N__4098\,
            I => \N__4092\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__4095\,
            I => \N__4086\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__4092\,
            I => \N__4086\
        );

    \I__542\ : InMux
    port map (
            O => \N__4091\,
            I => \N__4083\
        );

    \I__541\ : Span12Mux_s4_v
    port map (
            O => \N__4086\,
            I => \N__4080\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__4083\,
            I => n680
        );

    \I__539\ : Odrv12
    port map (
            O => \N__4080\,
            I => n680
        );

    \I__538\ : InMux
    port map (
            O => \N__4075\,
            I => \N__4071\
        );

    \I__537\ : InMux
    port map (
            O => \N__4074\,
            I => \N__4068\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__4071\,
            I => \N__4065\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__4068\,
            I => \N__4062\
        );

    \I__534\ : Odrv4
    port map (
            O => \N__4065\,
            I => data_reg_0
        );

    \I__533\ : Odrv4
    port map (
            O => \N__4062\,
            I => data_reg_0
        );

    \I__532\ : IoInMux
    port map (
            O => \N__4057\,
            I => \N__4054\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__4054\,
            I => \N__4051\
        );

    \I__530\ : Span4Mux_s3_v
    port map (
            O => \N__4051\,
            I => \N__4048\
        );

    \I__529\ : Odrv4
    port map (
            O => \N__4048\,
            I => output_axis_tdata_c_0
        );

    \I__528\ : InMux
    port map (
            O => \N__4045\,
            I => \N__4042\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__4042\,
            I => \N__4039\
        );

    \I__526\ : Span4Mux_v
    port map (
            O => \N__4039\,
            I => \N__4036\
        );

    \I__525\ : Odrv4
    port map (
            O => \N__4036\,
            I => rxd_c
        );

    \I__524\ : CascadeMux
    port map (
            O => \N__4033\,
            I => \uart_tx_inst.n910_cascade_\
        );

    \I__523\ : CascadeMux
    port map (
            O => \N__4030\,
            I => \N__4024\
        );

    \I__522\ : InMux
    port map (
            O => \N__4029\,
            I => \N__4019\
        );

    \I__521\ : InMux
    port map (
            O => \N__4028\,
            I => \N__4019\
        );

    \I__520\ : InMux
    port map (
            O => \N__4027\,
            I => \N__4016\
        );

    \I__519\ : InMux
    port map (
            O => \N__4024\,
            I => \N__4013\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__4019\,
            I => \uart_rx_inst.output_axis_tvalid_N_174\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__4016\,
            I => \uart_rx_inst.output_axis_tvalid_N_174\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__4013\,
            I => \uart_rx_inst.output_axis_tvalid_N_174\
        );

    \I__515\ : CascadeMux
    port map (
            O => \N__4006\,
            I => \n1711_cascade_\
        );

    \I__514\ : CascadeMux
    port map (
            O => \N__4003\,
            I => \n1220_cascade_\
        );

    \I__513\ : InMux
    port map (
            O => \N__4000\,
            I => \N__3994\
        );

    \I__512\ : InMux
    port map (
            O => \N__3999\,
            I => \N__3989\
        );

    \I__511\ : InMux
    port map (
            O => \N__3998\,
            I => \N__3989\
        );

    \I__510\ : InMux
    port map (
            O => \N__3997\,
            I => \N__3986\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__3994\,
            I => \uart_rx_inst.bit_cnt_3\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__3989\,
            I => \uart_rx_inst.bit_cnt_3\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__3986\,
            I => \uart_rx_inst.bit_cnt_3\
        );

    \I__506\ : CascadeMux
    port map (
            O => \N__3979\,
            I => \uart_rx_inst.output_axis_tvalid_N_172_cascade_\
        );

    \I__505\ : CascadeMux
    port map (
            O => \N__3976\,
            I => \uart_rx_inst.n232_cascade_\
        );

    \I__504\ : InMux
    port map (
            O => \N__3973\,
            I => \N__3969\
        );

    \I__503\ : InMux
    port map (
            O => \N__3972\,
            I => \N__3966\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__3969\,
            I => \N__3961\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__3966\,
            I => \N__3961\
        );

    \I__500\ : Span4Mux_v
    port map (
            O => \N__3961\,
            I => \N__3957\
        );

    \I__499\ : InMux
    port map (
            O => \N__3960\,
            I => \N__3954\
        );

    \I__498\ : Odrv4
    port map (
            O => \N__3957\,
            I => \uart_rx_inst.n1468\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__3954\,
            I => \uart_rx_inst.n1468\
        );

    \I__496\ : InMux
    port map (
            O => \N__3949\,
            I => \N__3946\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__3946\,
            I => \uart_rx_inst.n1502\
        );

    \I__494\ : InMux
    port map (
            O => \N__3943\,
            I => \N__3939\
        );

    \I__493\ : InMux
    port map (
            O => \N__3942\,
            I => \N__3936\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__3939\,
            I => \uart_rx_inst.n235\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__3936\,
            I => \uart_rx_inst.n235\
        );

    \I__490\ : CascadeMux
    port map (
            O => \N__3931\,
            I => \N__3927\
        );

    \I__489\ : InMux
    port map (
            O => \N__3930\,
            I => \N__3920\
        );

    \I__488\ : InMux
    port map (
            O => \N__3927\,
            I => \N__3917\
        );

    \I__487\ : InMux
    port map (
            O => \N__3926\,
            I => \N__3912\
        );

    \I__486\ : InMux
    port map (
            O => \N__3925\,
            I => \N__3912\
        );

    \I__485\ : InMux
    port map (
            O => \N__3924\,
            I => \N__3909\
        );

    \I__484\ : InMux
    port map (
            O => \N__3923\,
            I => \N__3906\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__3920\,
            I => \uart_rx_inst.bit_cnt_1\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__3917\,
            I => \uart_rx_inst.bit_cnt_1\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__3912\,
            I => \uart_rx_inst.bit_cnt_1\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__3909\,
            I => \uart_rx_inst.bit_cnt_1\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__3906\,
            I => \uart_rx_inst.bit_cnt_1\
        );

    \I__478\ : InMux
    port map (
            O => \N__3895\,
            I => \N__3888\
        );

    \I__477\ : InMux
    port map (
            O => \N__3894\,
            I => \N__3885\
        );

    \I__476\ : InMux
    port map (
            O => \N__3893\,
            I => \N__3880\
        );

    \I__475\ : InMux
    port map (
            O => \N__3892\,
            I => \N__3880\
        );

    \I__474\ : InMux
    port map (
            O => \N__3891\,
            I => \N__3877\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__3888\,
            I => \uart_rx_inst.bit_cnt_2\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__3885\,
            I => \uart_rx_inst.bit_cnt_2\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__3880\,
            I => \uart_rx_inst.bit_cnt_2\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__3877\,
            I => \uart_rx_inst.bit_cnt_2\
        );

    \I__469\ : CEMux
    port map (
            O => \N__3868\,
            I => \N__3864\
        );

    \I__468\ : CEMux
    port map (
            O => \N__3867\,
            I => \N__3861\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__3864\,
            I => \N__3858\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__3861\,
            I => \N__3855\
        );

    \I__465\ : Span4Mux_h
    port map (
            O => \N__3858\,
            I => \N__3851\
        );

    \I__464\ : Span4Mux_h
    port map (
            O => \N__3855\,
            I => \N__3848\
        );

    \I__463\ : InMux
    port map (
            O => \N__3854\,
            I => \N__3845\
        );

    \I__462\ : Odrv4
    port map (
            O => \N__3851\,
            I => n705
        );

    \I__461\ : Odrv4
    port map (
            O => \N__3848\,
            I => n705
        );

    \I__460\ : LocalMux
    port map (
            O => \N__3845\,
            I => n705
        );

    \I__459\ : CascadeMux
    port map (
            O => \N__3838\,
            I => \uart_rx_inst.n509_cascade_\
        );

    \I__458\ : InMux
    port map (
            O => \N__3835\,
            I => \N__3832\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__3832\,
            I => \uart_rx_inst.n31\
        );

    \I__456\ : InMux
    port map (
            O => \N__3829\,
            I => \N__3826\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__3826\,
            I => \uart_rx_inst.n33\
        );

    \I__454\ : CascadeMux
    port map (
            O => \N__3823\,
            I => \N__3800\
        );

    \I__453\ : InMux
    port map (
            O => \N__3822\,
            I => \N__3796\
        );

    \I__452\ : InMux
    port map (
            O => \N__3821\,
            I => \N__3779\
        );

    \I__451\ : InMux
    port map (
            O => \N__3820\,
            I => \N__3779\
        );

    \I__450\ : InMux
    port map (
            O => \N__3819\,
            I => \N__3779\
        );

    \I__449\ : InMux
    port map (
            O => \N__3818\,
            I => \N__3779\
        );

    \I__448\ : InMux
    port map (
            O => \N__3817\,
            I => \N__3779\
        );

    \I__447\ : InMux
    port map (
            O => \N__3816\,
            I => \N__3779\
        );

    \I__446\ : InMux
    port map (
            O => \N__3815\,
            I => \N__3779\
        );

    \I__445\ : InMux
    port map (
            O => \N__3814\,
            I => \N__3779\
        );

    \I__444\ : InMux
    port map (
            O => \N__3813\,
            I => \N__3766\
        );

    \I__443\ : InMux
    port map (
            O => \N__3812\,
            I => \N__3766\
        );

    \I__442\ : InMux
    port map (
            O => \N__3811\,
            I => \N__3766\
        );

    \I__441\ : InMux
    port map (
            O => \N__3810\,
            I => \N__3766\
        );

    \I__440\ : InMux
    port map (
            O => \N__3809\,
            I => \N__3766\
        );

    \I__439\ : InMux
    port map (
            O => \N__3808\,
            I => \N__3766\
        );

    \I__438\ : InMux
    port map (
            O => \N__3807\,
            I => \N__3761\
        );

    \I__437\ : InMux
    port map (
            O => \N__3806\,
            I => \N__3761\
        );

    \I__436\ : InMux
    port map (
            O => \N__3805\,
            I => \N__3750\
        );

    \I__435\ : InMux
    port map (
            O => \N__3804\,
            I => \N__3750\
        );

    \I__434\ : InMux
    port map (
            O => \N__3803\,
            I => \N__3750\
        );

    \I__433\ : InMux
    port map (
            O => \N__3800\,
            I => \N__3750\
        );

    \I__432\ : InMux
    port map (
            O => \N__3799\,
            I => \N__3750\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__3796\,
            I => \uart_rx_inst.n1479\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__3779\,
            I => \uart_rx_inst.n1479\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__3766\,
            I => \uart_rx_inst.n1479\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__3761\,
            I => \uart_rx_inst.n1479\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__3750\,
            I => \uart_rx_inst.n1479\
        );

    \I__426\ : CEMux
    port map (
            O => \N__3739\,
            I => \N__3735\
        );

    \I__425\ : CEMux
    port map (
            O => \N__3738\,
            I => \N__3730\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__3735\,
            I => \N__3727\
        );

    \I__423\ : CEMux
    port map (
            O => \N__3734\,
            I => \N__3724\
        );

    \I__422\ : CEMux
    port map (
            O => \N__3733\,
            I => \N__3721\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__3730\,
            I => \uart_rx_inst.n1045\
        );

    \I__420\ : Odrv4
    port map (
            O => \N__3727\,
            I => \uart_rx_inst.n1045\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__3724\,
            I => \uart_rx_inst.n1045\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__3721\,
            I => \uart_rx_inst.n1045\
        );

    \I__417\ : CascadeMux
    port map (
            O => \N__3712\,
            I => \uart_rx_inst.n30_cascade_\
        );

    \I__416\ : CascadeMux
    port map (
            O => \N__3709\,
            I => \uart_rx_inst.n32_cascade_\
        );

    \I__415\ : InMux
    port map (
            O => \N__3706\,
            I => \N__3703\
        );

    \I__414\ : LocalMux
    port map (
            O => \N__3703\,
            I => \uart_rx_inst.n34\
        );

    \I__413\ : CascadeMux
    port map (
            O => \N__3700\,
            I => \output_axis_tvalid_N_175_cascade_\
        );

    \I__412\ : CascadeMux
    port map (
            O => \N__3697\,
            I => \N__3691\
        );

    \I__411\ : CascadeMux
    port map (
            O => \N__3696\,
            I => \N__3686\
        );

    \I__410\ : CascadeMux
    port map (
            O => \N__3695\,
            I => \N__3683\
        );

    \I__409\ : InMux
    port map (
            O => \N__3694\,
            I => \N__3675\
        );

    \I__408\ : InMux
    port map (
            O => \N__3691\,
            I => \N__3675\
        );

    \I__407\ : InMux
    port map (
            O => \N__3690\,
            I => \N__3675\
        );

    \I__406\ : InMux
    port map (
            O => \N__3689\,
            I => \N__3666\
        );

    \I__405\ : InMux
    port map (
            O => \N__3686\,
            I => \N__3666\
        );

    \I__404\ : InMux
    port map (
            O => \N__3683\,
            I => \N__3666\
        );

    \I__403\ : InMux
    port map (
            O => \N__3682\,
            I => \N__3666\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__3675\,
            I => bit_cnt_2
        );

    \I__401\ : LocalMux
    port map (
            O => \N__3666\,
            I => bit_cnt_2
        );

    \I__400\ : InMux
    port map (
            O => \N__3661\,
            I => \N__3649\
        );

    \I__399\ : InMux
    port map (
            O => \N__3660\,
            I => \N__3649\
        );

    \I__398\ : InMux
    port map (
            O => \N__3659\,
            I => \N__3649\
        );

    \I__397\ : InMux
    port map (
            O => \N__3658\,
            I => \N__3642\
        );

    \I__396\ : InMux
    port map (
            O => \N__3657\,
            I => \N__3642\
        );

    \I__395\ : InMux
    port map (
            O => \N__3656\,
            I => \N__3642\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__3649\,
            I => \uart_tx_inst.bit_cnt_3\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__3642\,
            I => \uart_tx_inst.bit_cnt_3\
        );

    \I__392\ : CascadeMux
    port map (
            O => \N__3637\,
            I => \uart_tx_inst.n1723_cascade_\
        );

    \I__391\ : SRMux
    port map (
            O => \N__3634\,
            I => \N__3631\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__3631\,
            I => \N__3628\
        );

    \I__389\ : Odrv4
    port map (
            O => \N__3628\,
            I => \uart_rx_inst.n681\
        );

    \I__388\ : InMux
    port map (
            O => \N__3625\,
            I => \N__3622\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__3622\,
            I => \uart_tx_inst.n13\
        );

    \I__386\ : InMux
    port map (
            O => \N__3619\,
            I => \N__3616\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__3616\,
            I => \N__3613\
        );

    \I__384\ : Span4Mux_h
    port map (
            O => \N__3613\,
            I => \N__3610\
        );

    \I__383\ : Odrv4
    port map (
            O => \N__3610\,
            I => output_axis_tready_c
        );

    \I__382\ : IoInMux
    port map (
            O => \N__3607\,
            I => \N__3604\
        );

    \I__381\ : LocalMux
    port map (
            O => \N__3604\,
            I => \N__3601\
        );

    \I__380\ : Span4Mux_s3_v
    port map (
            O => \N__3601\,
            I => \N__3596\
        );

    \I__379\ : InMux
    port map (
            O => \N__3600\,
            I => \N__3593\
        );

    \I__378\ : InMux
    port map (
            O => \N__3599\,
            I => \N__3590\
        );

    \I__377\ : Odrv4
    port map (
            O => \N__3596\,
            I => output_axis_tvalid_c
        );

    \I__376\ : LocalMux
    port map (
            O => \N__3593\,
            I => output_axis_tvalid_c
        );

    \I__375\ : LocalMux
    port map (
            O => \N__3590\,
            I => output_axis_tvalid_c
        );

    \I__374\ : InMux
    port map (
            O => \N__3583\,
            I => \N__3579\
        );

    \I__373\ : InMux
    port map (
            O => \N__3582\,
            I => \N__3576\
        );

    \I__372\ : LocalMux
    port map (
            O => \N__3579\,
            I => \N__3573\
        );

    \I__371\ : LocalMux
    port map (
            O => \N__3576\,
            I => n1471
        );

    \I__370\ : Odrv4
    port map (
            O => \N__3573\,
            I => n1471
        );

    \I__369\ : CascadeMux
    port map (
            O => \N__3568\,
            I => \uart_tx_inst.n485_cascade_\
        );

    \I__368\ : CascadeMux
    port map (
            O => \N__3565\,
            I => \uart_tx_inst.n30_adj_196_cascade_\
        );

    \I__367\ : CascadeMux
    port map (
            O => \N__3562\,
            I => \uart_tx_inst.n34_cascade_\
        );

    \I__366\ : CascadeMux
    port map (
            O => \N__3559\,
            I => \uart_tx_inst.n189_cascade_\
        );

    \I__365\ : InMux
    port map (
            O => \N__3556\,
            I => \N__3552\
        );

    \I__364\ : CascadeMux
    port map (
            O => \N__3555\,
            I => \N__3545\
        );

    \I__363\ : LocalMux
    port map (
            O => \N__3552\,
            I => \N__3542\
        );

    \I__362\ : InMux
    port map (
            O => \N__3551\,
            I => \N__3539\
        );

    \I__361\ : InMux
    port map (
            O => \N__3550\,
            I => \N__3536\
        );

    \I__360\ : InMux
    port map (
            O => \N__3549\,
            I => \N__3533\
        );

    \I__359\ : InMux
    port map (
            O => \N__3548\,
            I => \N__3528\
        );

    \I__358\ : InMux
    port map (
            O => \N__3545\,
            I => \N__3528\
        );

    \I__357\ : Odrv4
    port map (
            O => \N__3542\,
            I => \uart_tx_inst.bit_cnt_0\
        );

    \I__356\ : LocalMux
    port map (
            O => \N__3539\,
            I => \uart_tx_inst.bit_cnt_0\
        );

    \I__355\ : LocalMux
    port map (
            O => \N__3536\,
            I => \uart_tx_inst.bit_cnt_0\
        );

    \I__354\ : LocalMux
    port map (
            O => \N__3533\,
            I => \uart_tx_inst.bit_cnt_0\
        );

    \I__353\ : LocalMux
    port map (
            O => \N__3528\,
            I => \uart_tx_inst.bit_cnt_0\
        );

    \I__352\ : CascadeMux
    port map (
            O => \N__3517\,
            I => \N__3514\
        );

    \I__351\ : InMux
    port map (
            O => \N__3514\,
            I => \N__3511\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__3511\,
            I => \uart_tx_inst.n7_adj_195\
        );

    \I__349\ : InMux
    port map (
            O => \N__3508\,
            I => \N__3499\
        );

    \I__348\ : InMux
    port map (
            O => \N__3507\,
            I => \N__3494\
        );

    \I__347\ : InMux
    port map (
            O => \N__3506\,
            I => \N__3494\
        );

    \I__346\ : InMux
    port map (
            O => \N__3505\,
            I => \N__3485\
        );

    \I__345\ : InMux
    port map (
            O => \N__3504\,
            I => \N__3485\
        );

    \I__344\ : InMux
    port map (
            O => \N__3503\,
            I => \N__3485\
        );

    \I__343\ : InMux
    port map (
            O => \N__3502\,
            I => \N__3485\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__3499\,
            I => \uart_tx_inst.bit_cnt_1\
        );

    \I__341\ : LocalMux
    port map (
            O => \N__3494\,
            I => \uart_tx_inst.bit_cnt_1\
        );

    \I__340\ : LocalMux
    port map (
            O => \N__3485\,
            I => \uart_tx_inst.bit_cnt_1\
        );

    \I__339\ : CascadeMux
    port map (
            O => \N__3478\,
            I => \uart_tx_inst.n15_cascade_\
        );

    \I__338\ : CascadeMux
    port map (
            O => \N__3475\,
            I => \n1167_cascade_\
        );

    \I__337\ : InMux
    port map (
            O => \N__3472\,
            I => \N__3469\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__3469\,
            I => n1698
        );

    \I__335\ : CascadeMux
    port map (
            O => \N__3466\,
            I => \uart_rx_inst.n677_cascade_\
        );

    \I__334\ : CascadeMux
    port map (
            O => \N__3463\,
            I => \uart_rx_inst.n607_cascade_\
        );

    \I__333\ : CascadeMux
    port map (
            O => \N__3460\,
            I => \uart_rx_inst.n603_cascade_\
        );

    \I__332\ : CEMux
    port map (
            O => \N__3457\,
            I => \N__3454\
        );

    \I__331\ : LocalMux
    port map (
            O => \N__3454\,
            I => \N__3451\
        );

    \I__330\ : Odrv12
    port map (
            O => \N__3451\,
            I => \uart_rx_inst.n984\
        );

    \I__329\ : CascadeMux
    port map (
            O => \N__3448\,
            I => \n705_cascade_\
        );

    \I__328\ : CascadeMux
    port map (
            O => \N__3445\,
            I => \uart_tx_inst.n7_cascade_\
        );

    \I__327\ : SRMux
    port map (
            O => \N__3442\,
            I => \N__3439\
        );

    \I__326\ : LocalMux
    port map (
            O => \N__3439\,
            I => \N__3436\
        );

    \I__325\ : Span4Mux_s0_v
    port map (
            O => \N__3436\,
            I => \N__3432\
        );

    \I__324\ : InMux
    port map (
            O => \N__3435\,
            I => \N__3429\
        );

    \I__323\ : Odrv4
    port map (
            O => \N__3432\,
            I => n1165
        );

    \I__322\ : LocalMux
    port map (
            O => \N__3429\,
            I => n1165
        );

    \I__321\ : CascadeMux
    port map (
            O => \N__3424\,
            I => \N__3421\
        );

    \I__320\ : InMux
    port map (
            O => \N__3421\,
            I => \N__3418\
        );

    \I__319\ : LocalMux
    port map (
            O => \N__3418\,
            I => n4
        );

    \I__318\ : InMux
    port map (
            O => \N__3415\,
            I => \N__3412\
        );

    \I__317\ : LocalMux
    port map (
            O => \N__3412\,
            I => \uart_tx_inst.n613\
        );

    \I__316\ : CEMux
    port map (
            O => \N__3409\,
            I => \N__3406\
        );

    \I__315\ : LocalMux
    port map (
            O => \N__3406\,
            I => \N__3402\
        );

    \I__314\ : CEMux
    port map (
            O => \N__3405\,
            I => \N__3399\
        );

    \I__313\ : Span4Mux_v
    port map (
            O => \N__3402\,
            I => \N__3394\
        );

    \I__312\ : LocalMux
    port map (
            O => \N__3399\,
            I => \N__3394\
        );

    \I__311\ : Span4Mux_s1_v
    port map (
            O => \N__3394\,
            I => \N__3390\
        );

    \I__310\ : InMux
    port map (
            O => \N__3393\,
            I => \N__3387\
        );

    \I__309\ : Odrv4
    port map (
            O => \N__3390\,
            I => n707
        );

    \I__308\ : LocalMux
    port map (
            O => \N__3387\,
            I => n707
        );

    \I__307\ : IoInMux
    port map (
            O => \N__3382\,
            I => \N__3379\
        );

    \I__306\ : LocalMux
    port map (
            O => \N__3379\,
            I => \N__3376\
        );

    \I__305\ : IoSpan4Mux
    port map (
            O => \N__3376\,
            I => \N__3373\
        );

    \I__304\ : Span4Mux_s0_v
    port map (
            O => \N__3373\,
            I => \N__3370\
        );

    \I__303\ : Odrv4
    port map (
            O => \N__3370\,
            I => rx_overrun_error_c
        );

    \I__302\ : CEMux
    port map (
            O => \N__3367\,
            I => \N__3364\
        );

    \I__301\ : LocalMux
    port map (
            O => \N__3364\,
            I => \N__3361\
        );

    \I__300\ : Odrv4
    port map (
            O => \N__3361\,
            I => \uart_tx_inst.n721\
        );

    \I__299\ : IoInMux
    port map (
            O => \N__3358\,
            I => \N__3355\
        );

    \I__298\ : LocalMux
    port map (
            O => \N__3355\,
            I => \N__3352\
        );

    \I__297\ : Span4Mux_s1_v
    port map (
            O => \N__3352\,
            I => \N__3348\
        );

    \I__296\ : InMux
    port map (
            O => \N__3351\,
            I => \N__3345\
        );

    \I__295\ : Odrv4
    port map (
            O => \N__3348\,
            I => input_axis_tready_c
        );

    \I__294\ : LocalMux
    port map (
            O => \N__3345\,
            I => input_axis_tready_c
        );

    \I__293\ : CEMux
    port map (
            O => \N__3340\,
            I => \N__3337\
        );

    \I__292\ : LocalMux
    port map (
            O => \N__3337\,
            I => \N__3334\
        );

    \I__291\ : Span4Mux_h
    port map (
            O => \N__3334\,
            I => \N__3331\
        );

    \I__290\ : Odrv4
    port map (
            O => \N__3331\,
            I => \uart_tx_inst.n701\
        );

    \I__289\ : SRMux
    port map (
            O => \N__3328\,
            I => \N__3325\
        );

    \I__288\ : LocalMux
    port map (
            O => \N__3325\,
            I => \uart_tx_inst.n535\
        );

    \I__287\ : IoInMux
    port map (
            O => \N__3322\,
            I => \N__3319\
        );

    \I__286\ : LocalMux
    port map (
            O => \N__3319\,
            I => \N__3316\
        );

    \I__285\ : Span12Mux_s5_v
    port map (
            O => \N__3316\,
            I => \N__3313\
        );

    \I__284\ : Odrv12
    port map (
            O => \N__3313\,
            I => rx_busy_c
        );

    \I__283\ : CascadeMux
    port map (
            O => \N__3310\,
            I => \n588_cascade_\
        );

    \I__282\ : CascadeMux
    port map (
            O => \N__3307\,
            I => \n707_cascade_\
        );

    \I__281\ : IoInMux
    port map (
            O => \N__3304\,
            I => \N__3301\
        );

    \I__280\ : LocalMux
    port map (
            O => \N__3301\,
            I => tx_busy_c
        );

    \IN_MUX_bfv_12_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_5_0_\
        );

    \IN_MUX_bfv_12_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \uart_tx_inst.n1589\,
            carryinitout => \bfn_12_6_0_\
        );

    \IN_MUX_bfv_11_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_2_0_\
        );

    \IN_MUX_bfv_11_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \uart_tx_inst.n1553\,
            carryinitout => \bfn_11_3_0_\
        );

    \IN_MUX_bfv_11_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \uart_tx_inst.n1561\,
            carryinitout => \bfn_11_4_0_\
        );

    \IN_MUX_bfv_9_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_5_0_\
        );

    \IN_MUX_bfv_9_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \uart_rx_inst.n1571\,
            carryinitout => \bfn_9_6_0_\
        );

    \IN_MUX_bfv_9_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \uart_rx_inst.n1579\,
            carryinitout => \bfn_9_7_0_\
        );

    \IN_MUX_bfv_11_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_5_0_\
        );

    \IN_MUX_bfv_11_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \uart_rx_inst.n1537\,
            carryinitout => \bfn_11_6_0_\
        );

    \IN_MUX_bfv_11_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \uart_rx_inst.n1545\,
            carryinitout => \bfn_11_7_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \uart_tx_inst.busy_reg_53_LC_5_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7660\,
            lcout => tx_busy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7365\,
            ce => \N__3367\,
            sr => \N__7188\
        );

    \uart_tx_inst.i1_2_lut_3_lut_LC_6_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__7185\,
            in1 => \N__7485\,
            in2 => \_gnd_net_\,
            in3 => \N__6708\,
            lcout => \uart_tx_inst.n701\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.i1_3_lut_adj_25_LC_6_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011101"
        )
    port map (
            in0 => \N__6709\,
            in1 => \N__7186\,
            in2 => \_gnd_net_\,
            in3 => \N__7486\,
            lcout => \uart_tx_inst.n721\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.i407_2_lut_LC_6_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__7187\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6707\,
            lcout => \uart_tx_inst.n535\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.input_axis_tready_reg_49_LC_6_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__7649\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3351\,
            lcout => input_axis_tready_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7366\,
            ce => \N__3340\,
            sr => \N__3328\
        );

    \uart_rx_inst.busy_reg_86_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5291\,
            lcout => rx_busy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7354\,
            ce => \N__3457\,
            sr => \N__7237\
        );

    \CONSTANT_ONE_LUT4_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.bit_cnt__i1_LC_7_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3556\,
            in2 => \_gnd_net_\,
            in3 => \N__3508\,
            lcout => \uart_tx_inst.bit_cnt_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7373\,
            ce => \N__3405\,
            sr => \N__3442\
        );

    \uart_tx_inst.i2_2_lut_4_lut_LC_7_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__3657\,
            in1 => \N__3503\,
            in2 => \N__3695\,
            in3 => \N__7430\,
            lcout => OPEN,
            ltout => \n588_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101110"
        )
    port map (
            in0 => \N__7161\,
            in1 => \N__3582\,
            in2 => \N__3310\,
            in3 => \N__6667\,
            lcout => n707,
            ltout => \n707_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.i1035_4_lut_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011010000"
        )
    port map (
            in0 => \N__7484\,
            in1 => \N__7162\,
            in2 => \N__3307\,
            in3 => \N__7431\,
            lcout => n1165,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.i1_2_lut_4_lut_adj_24_LC_7_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3502\,
            in1 => \N__3682\,
            in2 => \N__3555\,
            in3 => \N__3656\,
            lcout => \uart_tx_inst.n7\,
            ltout => \uart_tx_inst.n7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.i1343_2_lut_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3445\,
            in3 => \N__7645\,
            lcout => n1471,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.bit_cnt__i2_LC_7_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011000110"
        )
    port map (
            in0 => \N__3393\,
            in1 => \N__3689\,
            in2 => \N__3424\,
            in3 => \N__3435\,
            lcout => bit_cnt_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7370\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.i1_3_lut_4_lut_LC_7_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010110"
        )
    port map (
            in0 => \N__3658\,
            in1 => \N__3505\,
            in2 => \N__3696\,
            in3 => \N__3548\,
            lcout => \uart_tx_inst.n613\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.i266_2_lut_LC_7_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__3504\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3550\,
            lcout => n4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.bit_cnt__i3_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000111110000"
        )
    port map (
            in0 => \N__7437\,
            in1 => \N__3415\,
            in2 => \N__7659\,
            in3 => \N__7519\,
            lcout => \uart_tx_inst.bit_cnt_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7367\,
            ce => \N__3409\,
            sr => \N__7231\
        );

    \uart_tx_inst.bit_cnt__i0_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000001110100"
        )
    port map (
            in0 => \N__7436\,
            in1 => \N__7518\,
            in2 => \N__7658\,
            in3 => \N__3551\,
            lcout => \uart_tx_inst.bit_cnt_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7367\,
            ce => \N__3409\,
            sr => \N__7231\
        );

    \uart_rx_inst.overrun_error_reg_87_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3600\,
            lcout => rx_overrun_error_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7362\,
            ce => 'H',
            sr => \N__3634\
        );

    \uart_rx_inst.prescale_reg__i5_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__6181\,
            in1 => \N__3804\,
            in2 => \_gnd_net_\,
            in3 => \N__4384\,
            lcout => \uart_rx_inst.prescale_reg_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7359\,
            ce => \N__3733\,
            sr => \N__7239\
        );

    \uart_rx_inst.prescale_reg__i4_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__3803\,
            in1 => \N__5866\,
            in2 => \_gnd_net_\,
            in3 => \N__4423\,
            lcout => \uart_rx_inst.prescale_reg_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7359\,
            ce => \N__3733\,
            sr => \N__7239\
        );

    \uart_rx_inst.prescale_reg__i8_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__6142\,
            in1 => \N__3805\,
            in2 => \_gnd_net_\,
            in3 => \N__4774\,
            lcout => \uart_rx_inst.prescale_reg_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7359\,
            ce => \N__3733\,
            sr => \N__7239\
        );

    \uart_rx_inst.i1585_4_lut_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111011101"
        )
    port map (
            in0 => \N__4596\,
            in1 => \N__7243\,
            in2 => \N__3823\,
            in3 => \N__3972\,
            lcout => \uart_rx_inst.n1648\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i1011_2_lut_4_lut_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__7242\,
            in1 => \N__3799\,
            in2 => \_gnd_net_\,
            in3 => \N__4595\,
            lcout => \uart_rx_inst.n1141\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i1596_4_lut_4_lut_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011111111"
        )
    port map (
            in0 => \N__3973\,
            in1 => \N__3806\,
            in2 => \N__7263\,
            in3 => \N__4597\,
            lcout => \uart_rx_inst.n1045\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i854_2_lut_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__3807\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7236\,
            lcout => \uart_rx_inst.n984\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.prescale_reg__i2_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__5893\,
            in1 => \N__3822\,
            in2 => \_gnd_net_\,
            in3 => \N__4477\,
            lcout => \uart_rx_inst.prescale_reg_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7355\,
            ce => \N__3734\,
            sr => \N__7232\
        );

    \uart_rx_inst.i1568_2_lut_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6904\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6287\,
            lcout => \uart_rx_inst.n1756\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i1571_2_lut_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6288\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8002\,
            lcout => \uart_rx_inst.n1744\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__7252\,
            in1 => \N__3472\,
            in2 => \_gnd_net_\,
            in3 => \N__4127\,
            lcout => n705,
            ltout => \n705_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i1037_4_lut_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011110000"
        )
    port map (
            in0 => \N__7253\,
            in1 => \N__4027\,
            in2 => \N__3448\,
            in3 => \N__6311\,
            lcout => n1167,
            ltout => \n1167_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.bit_cnt__i0_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4257\,
            in2 => \N__3475\,
            in3 => \N__3854\,
            lcout => bit_cnt_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7352\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i1_4_lut_4_lut_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001011001110"
        )
    port map (
            in0 => \N__5293\,
            in1 => \N__4206\,
            in2 => \N__4270\,
            in3 => \N__3960\,
            lcout => n1698,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i2_3_lut_adj_22_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__4000\,
            in1 => \N__3894\,
            in2 => \_gnd_net_\,
            in3 => \N__3923\,
            lcout => \uart_rx_inst.n677\,
            ltout => \uart_rx_inst.n677_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i1_2_lut_adj_23_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3466\,
            in3 => \N__4253\,
            lcout => \uart_rx_inst.output_axis_tvalid_N_174\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i1_3_lut_4_lut_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010110"
        )
    port map (
            in0 => \N__3999\,
            in1 => \N__3893\,
            in2 => \N__3931\,
            in3 => \N__4263\,
            lcout => OPEN,
            ltout => \uart_rx_inst.n607_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.bit_cnt__i3_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100001011101"
        )
    port map (
            in0 => \N__4029\,
            in1 => \N__6313\,
            in2 => \N__3463\,
            in3 => \N__5296\,
            lcout => \uart_rx_inst.bit_cnt_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7356\,
            ce => \N__3867\,
            sr => \N__7264\
        );

    \uart_rx_inst.i1_2_lut_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4262\,
            in2 => \_gnd_net_\,
            in3 => \N__3926\,
            lcout => OPEN,
            ltout => \uart_rx_inst.n603_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.bit_cnt__i1_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100001011101"
        )
    port map (
            in0 => \N__4028\,
            in1 => \N__6312\,
            in2 => \N__3460\,
            in3 => \N__5295\,
            lcout => \uart_rx_inst.bit_cnt_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7356\,
            ce => \N__3867\,
            sr => \N__7264\
        );

    \uart_rx_inst.i209_2_lut_3_lut_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__3998\,
            in1 => \N__3892\,
            in2 => \_gnd_net_\,
            in3 => \N__3925\,
            lcout => \uart_rx_inst.output_axis_tvalid_N_173\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.i319_4_lut_LC_8_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101110"
        )
    port map (
            in0 => \N__6554\,
            in1 => \N__3583\,
            in2 => \N__3517\,
            in3 => \N__6668\,
            lcout => \uart_tx_inst.n485\,
            ltout => \uart_tx_inst.n485_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.i787_3_lut_LC_8_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8803\,
            in2 => \N__3568\,
            in3 => \N__6052\,
            lcout => \uart_tx_inst.n915\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.i11_4_lut_LC_8_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5850\,
            in1 => \N__5754\,
            in2 => \N__5928\,
            in3 => \N__5587\,
            lcout => OPEN,
            ltout => \uart_tx_inst.n30_adj_196_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.i15_4_lut_LC_8_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5724\,
            in1 => \N__5823\,
            in2 => \N__3565\,
            in3 => \N__6063\,
            lcout => OPEN,
            ltout => \uart_tx_inst.n34_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.i18_4_lut_LC_8_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4300\,
            in1 => \N__6196\,
            in2 => \N__3562\,
            in3 => \N__5374\,
            lcout => \input_axis_tready_N_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.i2_3_lut_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__7133\,
            in1 => \N__6569\,
            in2 => \_gnd_net_\,
            in3 => \N__6669\,
            lcout => \uart_tx_inst.n189\,
            ltout => \uart_tx_inst.n189_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.data_reg_i0_i8_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__7605\,
            in1 => \N__7563\,
            in2 => \N__3559\,
            in3 => \N__7483\,
            lcout => \uart_tx_inst.data_reg_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7375\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.i1_2_lut_4_lut_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__3660\,
            in1 => \N__3549\,
            in2 => \N__3697\,
            in3 => \N__3507\,
            lcout => \uart_tx_inst.n7_adj_195\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.i1_4_lut_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__3506\,
            in1 => \N__3690\,
            in2 => \_gnd_net_\,
            in3 => \N__3659\,
            lcout => \uart_tx_inst.n15\,
            ltout => \uart_tx_inst.n15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.i146_3_lut_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100001010"
        )
    port map (
            in0 => \N__7481\,
            in1 => \_gnd_net_\,
            in2 => \N__3478\,
            in3 => \N__7606\,
            lcout => \uart_tx_inst.n165\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.i1527_2_lut_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3694\,
            in2 => \_gnd_net_\,
            in3 => \N__3661\,
            lcout => OPEN,
            ltout => \uart_tx_inst.n1723_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.i29_4_lut_LC_8_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111011101110"
        )
    port map (
            in0 => \N__7482\,
            in1 => \N__7607\,
            in2 => \N__3637\,
            in3 => \N__7432\,
            lcout => \uart_tx_inst.n13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i1587_2_lut_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7176\,
            in2 => \_gnd_net_\,
            in3 => \N__4098\,
            lcout => \uart_rx_inst.n681\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.i1_3_lut_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__7177\,
            in1 => \N__3625\,
            in2 => \_gnd_net_\,
            in3 => \N__6721\,
            lcout => \uart_tx_inst.n719\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.output_axis_tvalid_reg_82_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__3619\,
            in1 => \N__3599\,
            in2 => \_gnd_net_\,
            in3 => \N__4099\,
            lcout => output_axis_tvalid_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7368\,
            ce => 'H',
            sr => \N__7163\
        );

    \uart_rx_inst.prescale_reg__i3_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__5878\,
            in1 => \N__3818\,
            in2 => \_gnd_net_\,
            in3 => \N__4450\,
            lcout => \uart_rx_inst.prescale_reg_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7363\,
            ce => \N__3739\,
            sr => \N__7241\
        );

    \uart_rx_inst.prescale_reg__i18_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__3817\,
            in1 => \N__6334\,
            in2 => \_gnd_net_\,
            in3 => \N__4834\,
            lcout => \uart_rx_inst.prescale_reg_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7363\,
            ce => \N__3739\,
            sr => \N__7241\
        );

    \uart_rx_inst.prescale_reg__i14_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__6397\,
            in1 => \N__3816\,
            in2 => \_gnd_net_\,
            in3 => \N__4606\,
            lcout => \uart_rx_inst.prescale_reg_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7363\,
            ce => \N__3739\,
            sr => \N__7241\
        );

    \uart_rx_inst.prescale_reg__i11_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__3815\,
            in1 => \N__6100\,
            in2 => \_gnd_net_\,
            in3 => \N__4678\,
            lcout => \uart_rx_inst.prescale_reg_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7363\,
            ce => \N__3739\,
            sr => \N__7241\
        );

    \uart_rx_inst.prescale_reg__i10_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__6115\,
            in1 => \N__3814\,
            in2 => \_gnd_net_\,
            in3 => \N__4702\,
            lcout => \uart_rx_inst.prescale_reg_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7363\,
            ce => \N__3739\,
            sr => \N__7241\
        );

    \uart_rx_inst.prescale_reg__i9_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__3821\,
            in1 => \N__6127\,
            in2 => \_gnd_net_\,
            in3 => \N__4738\,
            lcout => \uart_rx_inst.prescale_reg_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7363\,
            ce => \N__3739\,
            sr => \N__7241\
        );

    \uart_rx_inst.prescale_reg__i7_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__6154\,
            in1 => \N__3820\,
            in2 => \_gnd_net_\,
            in3 => \N__4336\,
            lcout => \uart_rx_inst.prescale_reg_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7363\,
            ce => \N__3739\,
            sr => \N__7241\
        );

    \uart_rx_inst.prescale_reg__i6_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__3819\,
            in1 => \_gnd_net_\,
            in2 => \N__6169\,
            in3 => \N__4357\,
            lcout => \uart_rx_inst.prescale_reg_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7363\,
            ce => \N__3739\,
            sr => \N__7241\
        );

    \uart_rx_inst.i1351_2_lut_3_lut_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__4273\,
            in1 => \N__4212\,
            in2 => \_gnd_net_\,
            in3 => \N__4125\,
            lcout => \uart_rx_inst.n1479\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i11_4_lut_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4848\,
            in1 => \N__4461\,
            in2 => \N__4717\,
            in3 => \N__4368\,
            lcout => OPEN,
            ltout => \uart_rx_inst.n30_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i15_4_lut_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4689\,
            in1 => \N__4347\,
            in2 => \N__3712\,
            in3 => \N__4617\,
            lcout => \uart_rx_inst.n34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i13_4_lut_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4575\,
            in1 => \N__4434\,
            in2 => \N__4791\,
            in3 => \N__4395\,
            lcout => OPEN,
            ltout => \uart_rx_inst.n32_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i18_4_lut_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3829\,
            in1 => \N__3835\,
            in2 => \N__3709\,
            in3 => \N__3706\,
            lcout => \output_axis_tvalid_N_175\,
            ltout => \output_axis_tvalid_N_175_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i362_3_lut_4_lut_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001110"
        )
    port map (
            in0 => \N__4272\,
            in1 => \N__5292\,
            in2 => \N__3700\,
            in3 => \N__4211\,
            lcout => \uart_rx_inst.n509\,
            ltout => \uart_rx_inst.n509_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i584_1_lut_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3838\,
            in3 => \_gnd_net_\,
            lcout => \uart_rx_inst.n712\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i12_4_lut_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4962\,
            in1 => \N__5013\,
            in2 => \N__4993\,
            in3 => \N__4641\,
            lcout => \uart_rx_inst.n31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.prescale_reg__i13_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__6412\,
            in1 => \N__3810\,
            in2 => \_gnd_net_\,
            in3 => \N__4630\,
            lcout => \uart_rx_inst.prescale_reg_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7357\,
            ce => \N__3738\,
            sr => \N__7244\
        );

    \uart_rx_inst.prescale_reg__i15_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__3811\,
            in1 => \N__6382\,
            in2 => \_gnd_net_\,
            in3 => \N__5002\,
            lcout => \uart_rx_inst.prescale_reg_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7357\,
            ce => \N__3738\,
            sr => \N__7244\
        );

    \uart_rx_inst.prescale_reg__i17_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__6352\,
            in1 => \N__3813\,
            in2 => \_gnd_net_\,
            in3 => \N__4951\,
            lcout => \uart_rx_inst.prescale_reg_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7357\,
            ce => \N__3738\,
            sr => \N__7244\
        );

    \uart_rx_inst.prescale_reg__i16_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__3812\,
            in1 => \N__6367\,
            in2 => \_gnd_net_\,
            in3 => \N__4978\,
            lcout => \uart_rx_inst.prescale_reg_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7357\,
            ce => \N__3738\,
            sr => \N__7244\
        );

    \uart_rx_inst.prescale_reg__i1_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3808\,
            in2 => \_gnd_net_\,
            in3 => \N__4510\,
            lcout => \uart_rx_inst.prescale_reg_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7357\,
            ce => \N__3738\,
            sr => \N__7244\
        );

    \uart_rx_inst.i14_4_lut_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4521\,
            in1 => \N__4488\,
            in2 => \N__4759\,
            in3 => \N__4668\,
            lcout => \uart_rx_inst.n33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.prescale_reg__i12_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3809\,
            in2 => \N__4657\,
            in3 => \N__6085\,
            lcout => \uart_rx_inst.prescale_reg_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7357\,
            ce => \N__3738\,
            sr => \N__7244\
        );

    \uart_rx_inst.i1516_4_lut_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101011100"
        )
    port map (
            in0 => \N__3942\,
            in1 => \N__5271\,
            in2 => \N__4030\,
            in3 => \N__3949\,
            lcout => n1711,
            ltout => \n1711_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i1384_3_lut_4_lut_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111000"
        )
    port map (
            in0 => \N__3943\,
            in1 => \N__4261\,
            in2 => \N__4006\,
            in3 => \N__4210\,
            lcout => n1220,
            ltout => \n1220_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.data_reg__i7_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000010000000"
        )
    port map (
            in0 => \N__5111\,
            in1 => \N__5355\,
            in2 => \N__4003\,
            in3 => \N__5272\,
            lcout => data_reg_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7353\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i208_2_lut_3_lut_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__3997\,
            in1 => \N__3891\,
            in2 => \_gnd_net_\,
            in3 => \N__3924\,
            lcout => \uart_rx_inst.output_axis_tvalid_N_172\,
            ltout => \uart_rx_inst.output_axis_tvalid_N_172_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i149_3_lut_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011111010"
        )
    port map (
            in0 => \N__4159\,
            in1 => \_gnd_net_\,
            in2 => \N__3979\,
            in3 => \N__5269\,
            lcout => \uart_rx_inst.n232\,
            ltout => \uart_rx_inst.n232_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i1340_3_lut_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011110000"
        )
    port map (
            in0 => \N__5270\,
            in1 => \_gnd_net_\,
            in2 => \N__3976\,
            in3 => \N__4160\,
            lcout => \uart_rx_inst.n1468\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i1374_2_lut_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__7245\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4126\,
            lcout => \uart_rx_inst.n1502\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i78_2_lut_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4173\,
            in2 => \_gnd_net_\,
            in3 => \N__4161\,
            lcout => \uart_rx_inst.n235\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.bit_cnt__i2_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010011001"
        )
    port map (
            in0 => \N__4264\,
            in1 => \N__3895\,
            in2 => \_gnd_net_\,
            in3 => \N__3930\,
            lcout => \uart_rx_inst.bit_cnt_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7358\,
            ce => \N__3868\,
            sr => \N__4285\
        );

    \uart_rx_inst.i2_4_lut_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__4271\,
            in1 => \N__4213\,
            in2 => \N__4180\,
            in3 => \N__4162\,
            lcout => n695,
            ltout => \n695_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.i1589_2_lut_3_lut_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101111"
        )
    port map (
            in0 => \N__7238\,
            in1 => \_gnd_net_\,
            in2 => \N__4144\,
            in3 => \N__4135\,
            lcout => n697,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.data_reg__i0_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__4074\,
            in1 => \N__5365\,
            in2 => \N__5494\,
            in3 => \N__5326\,
            lcout => data_reg_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7360\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i2_3_lut_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__4141\,
            in1 => \N__5282\,
            in2 => \_gnd_net_\,
            in3 => \N__4134\,
            lcout => n680,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__7255\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4091\,
            lcout => n703,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.output_axis_tdata_reg__i1_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4075\,
            lcout => output_axis_tdata_c_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7371\,
            ce => \N__5418\,
            sr => \N__7266\
        );

    \uart_rx_inst.rxd_reg_83_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4045\,
            lcout => rxd_reg,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7374\,
            ce => 'H',
            sr => \N__7267\
        );

    \uart_tx_inst.i782_3_lut_LC_9_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7714\,
            in1 => \N__5647\,
            in2 => \_gnd_net_\,
            in3 => \N__6775\,
            lcout => OPEN,
            ltout => \uart_tx_inst.n910_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.prescale_reg__i13_LC_9_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__6566\,
            in1 => \N__7784\,
            in2 => \N__4033\,
            in3 => \N__6690\,
            lcout => \uart_tx_inst.prescale_reg_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7379\,
            ce => \N__6476\,
            sr => \N__7072\
        );

    \uart_tx_inst.i792_3_lut_LC_9_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8701\,
            in1 => \N__6016\,
            in2 => \_gnd_net_\,
            in3 => \N__6776\,
            lcout => OPEN,
            ltout => \uart_tx_inst.n920_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.prescale_reg__i15_LC_9_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__6567\,
            in1 => \N__8775\,
            in2 => \N__4306\,
            in3 => \N__6691\,
            lcout => \uart_tx_inst.prescale_reg_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7379\,
            ce => \N__6476\,
            sr => \N__7072\
        );

    \uart_tx_inst.i802_3_lut_LC_9_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8491\,
            in1 => \N__5944\,
            in2 => \_gnd_net_\,
            in3 => \N__6777\,
            lcout => OPEN,
            ltout => \uart_tx_inst.n930_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.prescale_reg__i17_LC_9_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__6568\,
            in1 => \N__8571\,
            in2 => \N__4303\,
            in3 => \N__6692\,
            lcout => \uart_tx_inst.prescale_reg_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7379\,
            ce => \N__6476\,
            sr => \N__7072\
        );

    \uart_tx_inst.i12_4_lut_LC_9_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5955\,
            in1 => \N__6027\,
            in2 => \N__6000\,
            in3 => \N__5658\,
            lcout => \uart_tx_inst.n31_adj_199\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.i2_3_lut_4_lut_LC_9_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__6774\,
            in1 => \N__7073\,
            in2 => \N__6592\,
            in3 => \N__6689\,
            lcout => \uart_tx_inst.n873\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.prescale_reg__i14_LC_9_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__6570\,
            in1 => \N__4294\,
            in2 => \N__8872\,
            in3 => \N__6697\,
            lcout => \uart_tx_inst.prescale_reg_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7378\,
            ce => \N__6464\,
            sr => \N__7175\
        );

    \uart_tx_inst.i747_3_lut_LC_9_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8107\,
            in1 => \N__5836\,
            in2 => \_gnd_net_\,
            in3 => \N__6804\,
            lcout => OPEN,
            ltout => \uart_tx_inst.n875_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.prescale_reg__i6_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__8871\,
            in1 => \N__6574\,
            in2 => \N__4288\,
            in3 => \N__6698\,
            lcout => \uart_tx_inst.prescale_reg_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7378\,
            ce => \N__6464\,
            sr => \N__7175\
        );

    \uart_tx_inst.i752_3_lut_LC_9_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8080\,
            in1 => \N__5809\,
            in2 => \_gnd_net_\,
            in3 => \N__6805\,
            lcout => OPEN,
            ltout => \uart_tx_inst.n880_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.prescale_reg__i7_LC_9_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__8776\,
            in1 => \N__6575\,
            in2 => \N__4327\,
            in3 => \N__6699\,
            lcout => \uart_tx_inst.prescale_reg_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7378\,
            ce => \N__6464\,
            sr => \N__7175\
        );

    \uart_tx_inst.i767_3_lut_LC_9_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5743\,
            in1 => \N__7998\,
            in2 => \_gnd_net_\,
            in3 => \N__6806\,
            lcout => OPEN,
            ltout => \uart_tx_inst.n895_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.prescale_reg__i10_LC_9_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__8462\,
            in1 => \N__6573\,
            in2 => \N__4324\,
            in3 => \N__6696\,
            lcout => \uart_tx_inst.prescale_reg_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7378\,
            ce => \N__6464\,
            sr => \N__7175\
        );

    \uart_tx_inst.prescale_reg__i16_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__6571\,
            in1 => \N__4318\,
            in2 => \N__8674\,
            in3 => \N__6723\,
            lcout => \uart_tx_inst.prescale_reg_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7377\,
            ce => \N__6465\,
            sr => \N__7132\
        );

    \uart_tx_inst.prescale_reg__i18_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__6572\,
            in1 => \N__4312\,
            in2 => \N__8464\,
            in3 => \N__6724\,
            lcout => \uart_tx_inst.prescale_reg_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7377\,
            ce => \N__6465\,
            sr => \N__7132\
        );

    \uart_tx_inst.i772_3_lut_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7909\,
            in1 => \N__5707\,
            in2 => \_gnd_net_\,
            in3 => \N__6835\,
            lcout => OPEN,
            ltout => \uart_tx_inst.n900_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.prescale_reg__i11_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__7969\,
            in1 => \N__6576\,
            in2 => \N__4321\,
            in3 => \N__6722\,
            lcout => \uart_tx_inst.prescale_reg_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7377\,
            ce => \N__6465\,
            sr => \N__7132\
        );

    \uart_tx_inst.i797_3_lut_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8596\,
            in1 => \N__5977\,
            in2 => \_gnd_net_\,
            in3 => \N__6834\,
            lcout => \uart_tx_inst.n925\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.i807_3_lut_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6833\,
            in1 => \N__8131\,
            in2 => \_gnd_net_\,
            in3 => \N__5902\,
            lcout => \uart_tx_inst.n935\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.prescale_reg__i0_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__6322\,
            in1 => \N__4594\,
            in2 => \N__4576\,
            in3 => \N__4558\,
            lcout => \uart_rx_inst.prescale_reg_0\,
            ltout => OPEN,
            carryin => \bfn_9_5_0_\,
            carryout => \uart_rx_inst.n1564\,
            clk => \N__7369\,
            ce => \N__4555\,
            sr => \N__4543\
        );

    \uart_rx_inst.sub_10_add_2_3_lut_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__6320\,
            in1 => \N__4528\,
            in2 => \N__4934\,
            in3 => \N__4501\,
            lcout => \uart_rx_inst.n819\,
            ltout => OPEN,
            carryin => \uart_rx_inst.n1564\,
            carryout => \uart_rx_inst.n1565\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.sub_10_add_2_4_lut_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__6321\,
            in1 => \N__4901\,
            in2 => \N__4498\,
            in3 => \N__4465\,
            lcout => \uart_rx_inst.n814\,
            ltout => OPEN,
            carryin => \uart_rx_inst.n1565\,
            carryout => \uart_rx_inst.n1566\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.sub_10_add_2_5_lut_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__5050\,
            in1 => \N__4462\,
            in2 => \N__4935\,
            in3 => \N__4444\,
            lcout => \uart_rx_inst.n809\,
            ltout => OPEN,
            carryin => \uart_rx_inst.n1566\,
            carryout => \uart_rx_inst.n1567\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.sub_10_add_2_6_lut_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__5026\,
            in1 => \N__4905\,
            in2 => \N__4441\,
            in3 => \N__4414\,
            lcout => \uart_rx_inst.n804\,
            ltout => OPEN,
            carryin => \uart_rx_inst.n1567\,
            carryout => \uart_rx_inst.n1568\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.sub_10_add_2_7_lut_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__4411\,
            in1 => \N__4399\,
            in2 => \N__4936\,
            in3 => \N__4375\,
            lcout => \uart_rx_inst.n799\,
            ltout => OPEN,
            carryin => \uart_rx_inst.n1568\,
            carryout => \uart_rx_inst.n1569\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.sub_10_add_2_8_lut_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__5077\,
            in1 => \N__4909\,
            in2 => \N__4372\,
            in3 => \N__4351\,
            lcout => \uart_rx_inst.n794\,
            ltout => OPEN,
            carryin => \uart_rx_inst.n1569\,
            carryout => \uart_rx_inst.n1570\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.sub_10_add_2_9_lut_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__5035\,
            in1 => \N__4348\,
            in2 => \N__4937\,
            in3 => \N__4330\,
            lcout => \uart_rx_inst.n789\,
            ltout => OPEN,
            carryin => \uart_rx_inst.n1570\,
            carryout => \uart_rx_inst.n1571\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.sub_10_add_2_10_lut_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__4813\,
            in1 => \N__4795\,
            in2 => \N__4938\,
            in3 => \N__4762\,
            lcout => \uart_rx_inst.n784\,
            ltout => OPEN,
            carryin => \bfn_9_6_0_\,
            carryout => \uart_rx_inst.n1572\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.sub_10_add_2_11_lut_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__4825\,
            in1 => \N__4916\,
            in2 => \N__4758\,
            in3 => \N__4732\,
            lcout => \uart_rx_inst.n779\,
            ltout => OPEN,
            carryin => \uart_rx_inst.n1572\,
            carryout => \uart_rx_inst.n1573\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.sub_10_add_2_12_lut_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__4729\,
            in1 => \N__4716\,
            in2 => \N__4939\,
            in3 => \N__4696\,
            lcout => \uart_rx_inst.n774\,
            ltout => OPEN,
            carryin => \uart_rx_inst.n1573\,
            carryout => \uart_rx_inst.n1574\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.sub_10_add_2_13_lut_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__4801\,
            in1 => \N__4920\,
            in2 => \N__4693\,
            in3 => \N__4672\,
            lcout => \uart_rx_inst.n769\,
            ltout => OPEN,
            carryin => \uart_rx_inst.n1574\,
            carryout => \uart_rx_inst.n1575\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.sub_10_add_2_14_lut_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__6220\,
            in1 => \N__4669\,
            in2 => \N__4940\,
            in3 => \N__4648\,
            lcout => \uart_rx_inst.n764\,
            ltout => OPEN,
            carryin => \uart_rx_inst.n1575\,
            carryout => \uart_rx_inst.n1576\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.sub_10_add_2_15_lut_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__4807\,
            in1 => \N__4924\,
            in2 => \N__4645\,
            in3 => \N__4624\,
            lcout => \uart_rx_inst.n759\,
            ltout => OPEN,
            carryin => \uart_rx_inst.n1576\,
            carryout => \uart_rx_inst.n1577\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.sub_10_add_2_16_lut_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__5086\,
            in1 => \N__4621\,
            in2 => \N__4941\,
            in3 => \N__4600\,
            lcout => \uart_rx_inst.n754\,
            ltout => OPEN,
            carryin => \uart_rx_inst.n1577\,
            carryout => \uart_rx_inst.n1578\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.sub_10_add_2_17_lut_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__4819\,
            in1 => \N__4928\,
            in2 => \N__5017\,
            in3 => \N__4996\,
            lcout => \uart_rx_inst.n749\,
            ltout => OPEN,
            carryin => \uart_rx_inst.n1578\,
            carryout => \uart_rx_inst.n1579\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.sub_10_add_2_18_lut_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__5041\,
            in1 => \N__4992\,
            in2 => \N__4942\,
            in3 => \N__4972\,
            lcout => \uart_rx_inst.n744\,
            ltout => OPEN,
            carryin => \bfn_9_7_0_\,
            carryout => \uart_rx_inst.n1580\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.sub_10_add_2_19_lut_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__5059\,
            in1 => \N__4932\,
            in2 => \N__4969\,
            in3 => \N__4945\,
            lcout => \uart_rx_inst.n739\,
            ltout => OPEN,
            carryin => \uart_rx_inst.n1580\,
            carryout => \uart_rx_inst.n1581\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.sub_10_add_2_20_lut_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001110010"
        )
    port map (
            in0 => \N__4933\,
            in1 => \N__4852\,
            in2 => \N__5068\,
            in3 => \N__4837\,
            lcout => \uart_rx_inst.n729\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i1578_2_lut_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6302\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8028\,
            lcout => \uart_rx_inst.n1743\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i1569_2_lut_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8697\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6303\,
            lcout => \uart_rx_inst.n1740\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i1577_2_lut_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6300\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8056\,
            lcout => \uart_rx_inst.n1741\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i1574_2_lut_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7707\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6304\,
            lcout => \uart_rx_inst.n1747\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i1572_2_lut_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6301\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7905\,
            lcout => \uart_rx_inst.n1745\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i1563_2_lut_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8799\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6296\,
            lcout => \uart_rx_inst.n1750\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i1580_2_lut_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6295\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8106\,
            lcout => \uart_rx_inst.n1755\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i1565_2_lut_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8130\,
            in2 => \_gnd_net_\,
            in3 => \N__6298\,
            lcout => \uart_rx_inst.n1754\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i1576_2_lut_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6294\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8487\,
            lcout => \uart_rx_inst.n1751\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i1566_2_lut_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6961\,
            in2 => \_gnd_net_\,
            in3 => \N__6297\,
            lcout => \uart_rx_inst.n1758\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i1570_2_lut_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6299\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8595\,
            lcout => \uart_rx_inst.n1742\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i1581_2_lut_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8079\,
            in2 => \_gnd_net_\,
            in3 => \N__6293\,
            lcout => \uart_rx_inst.n1739\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i1567_2_lut_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6292\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6934\,
            lcout => \uart_rx_inst.n1757\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.data_reg__i2_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__5321\,
            in1 => \N__5453\,
            in2 => \N__5163\,
            in3 => \N__5362\,
            lcout => data_reg_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7361\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.data_reg__i5_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__5519\,
            in1 => \N__5361\,
            in2 => \N__5193\,
            in3 => \N__5324\,
            lcout => data_reg_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7361\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.data_reg__i3_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__5322\,
            in1 => \N__5553\,
            in2 => \N__5455\,
            in3 => \N__5363\,
            lcout => data_reg_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7361\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.data_reg__i1_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__5483\,
            in1 => \N__5359\,
            in2 => \N__5164\,
            in3 => \N__5320\,
            lcout => data_reg_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7361\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.data_reg__i6_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__5325\,
            in1 => \N__5186\,
            in2 => \N__5118\,
            in3 => \N__5364\,
            lcout => data_reg_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7361\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.data_reg__i4_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__5552\,
            in1 => \N__5360\,
            in2 => \N__5526\,
            in3 => \N__5323\,
            lcout => data_reg_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7361\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.frame_error_reg_88_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5294\,
            lcout => rx_frame_error_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7364\,
            ce => 'H',
            sr => \N__5206\
        );

    \uart_rx_inst.output_axis_tdata_reg__i7_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5194\,
            lcout => output_axis_tdata_c_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7372\,
            ce => \N__5408\,
            sr => \N__7254\
        );

    \uart_rx_inst.output_axis_tdata_reg__i3_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5162\,
            lcout => output_axis_tdata_c_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7372\,
            ce => \N__5408\,
            sr => \N__7254\
        );

    \uart_rx_inst.output_axis_tdata_reg__i8_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5122\,
            lcout => output_axis_tdata_c_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7372\,
            ce => \N__5408\,
            sr => \N__7254\
        );

    \uart_rx_inst.output_axis_tdata_reg__i5_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5557\,
            lcout => output_axis_tdata_c_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7372\,
            ce => \N__5408\,
            sr => \N__7254\
        );

    \uart_rx_inst.output_axis_tdata_reg__i6_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5527\,
            lcout => output_axis_tdata_c_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7372\,
            ce => \N__5408\,
            sr => \N__7254\
        );

    \uart_rx_inst.output_axis_tdata_reg__i2_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5493\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => output_axis_tdata_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7376\,
            ce => \N__5419\,
            sr => \N__7265\
        );

    \uart_rx_inst.output_axis_tdata_reg__i4_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5454\,
            lcout => output_axis_tdata_c_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7376\,
            ce => \N__5419\,
            sr => \N__7265\
        );

    \uart_tx_inst.i777_3_lut_LC_11_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6809\,
            in1 => \N__7813\,
            in2 => \_gnd_net_\,
            in3 => \N__5680\,
            lcout => OPEN,
            ltout => \uart_tx_inst.n905_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.prescale_reg__i12_LC_11_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__6594\,
            in1 => \N__7883\,
            in2 => \N__5380\,
            in3 => \N__6711\,
            lcout => \uart_tx_inst.prescale_reg_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7382\,
            ce => \N__6477\,
            sr => \N__7181\
        );

    \uart_tx_inst.i762_3_lut_LC_11_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6808\,
            in1 => \N__8029\,
            in2 => \_gnd_net_\,
            in3 => \N__5773\,
            lcout => OPEN,
            ltout => \uart_tx_inst.n890_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.prescale_reg__i9_LC_11_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__6595\,
            in1 => \N__8570\,
            in2 => \N__5377\,
            in3 => \N__6713\,
            lcout => \uart_tx_inst.prescale_reg_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7382\,
            ce => \N__6477\,
            sr => \N__7181\
        );

    \uart_tx_inst.i14_4_lut_LC_11_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5625\,
            in1 => \N__5610\,
            in2 => \N__5790\,
            in3 => \N__5691\,
            lcout => \uart_tx_inst.n33_adj_198\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.i732_3_lut_LC_11_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5572\,
            in1 => \N__6960\,
            in2 => \_gnd_net_\,
            in3 => \N__6810\,
            lcout => OPEN,
            ltout => \uart_tx_inst.n860_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.prescale_reg__i3_LC_11_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__6712\,
            in1 => \N__7970\,
            in2 => \N__5632\,
            in3 => \N__6596\,
            lcout => \uart_tx_inst.prescale_reg_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7382\,
            ce => \N__6477\,
            sr => \N__7181\
        );

    \uart_tx_inst.i1524_3_lut_4_lut_LC_11_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__6593\,
            in1 => \N__6807\,
            in2 => \N__7240\,
            in3 => \N__6710\,
            lcout => \uart_tx_inst.n1170\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.prescale_reg__i0_LC_11_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__6837\,
            in1 => \N__6208\,
            in2 => \_gnd_net_\,
            in3 => \N__5629\,
            lcout => \uart_tx_inst.prescale_reg_0\,
            ltout => OPEN,
            carryin => \bfn_11_2_0_\,
            carryout => \uart_tx_inst.n1546\,
            clk => \N__7380\,
            ce => \N__6481\,
            sr => \N__5596\
        );

    \uart_tx_inst.prescale_reg__i1_LC_11_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__6836\,
            in1 => \N__5626\,
            in2 => \N__8380\,
            in3 => \N__5614\,
            lcout => \uart_tx_inst.prescale_reg_1\,
            ltout => OPEN,
            carryin => \uart_tx_inst.n1546\,
            carryout => \uart_tx_inst.n1547\,
            clk => \N__7380\,
            ce => \N__6481\,
            sr => \N__5596\
        );

    \uart_tx_inst.prescale_reg__i2_LC_11_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__6838\,
            in1 => \N__5611\,
            in2 => \N__8374\,
            in3 => \N__5599\,
            lcout => \uart_tx_inst.prescale_reg_2\,
            ltout => OPEN,
            carryin => \uart_tx_inst.n1547\,
            carryout => \uart_tx_inst.n1548\,
            clk => \N__7380\,
            ce => \N__6481\,
            sr => \N__5596\
        );

    \uart_tx_inst.sub_5_add_2_5_lut_LC_11_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5586\,
            in2 => \N__8381\,
            in3 => \N__5566\,
            lcout => \uart_tx_inst.n33\,
            ltout => OPEN,
            carryin => \uart_tx_inst.n1548\,
            carryout => \uart_tx_inst.n1549\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.sub_5_add_2_6_lut_LC_11_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8366\,
            in2 => \N__6877\,
            in3 => \N__5563\,
            lcout => \uart_tx_inst.n32\,
            ltout => OPEN,
            carryin => \uart_tx_inst.n1549\,
            carryout => \uart_tx_inst.n1550\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.sub_5_add_2_7_lut_LC_11_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6850\,
            in2 => \N__8382\,
            in3 => \N__5560\,
            lcout => \uart_tx_inst.n31\,
            ltout => OPEN,
            carryin => \uart_tx_inst.n1550\,
            carryout => \uart_tx_inst.n1551\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.sub_5_add_2_8_lut_LC_11_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8370\,
            in2 => \N__5854\,
            in3 => \N__5827\,
            lcout => \uart_tx_inst.n30\,
            ltout => OPEN,
            carryin => \uart_tx_inst.n1551\,
            carryout => \uart_tx_inst.n1552\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.sub_5_add_2_9_lut_LC_11_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5824\,
            in2 => \N__8383\,
            in3 => \N__5800\,
            lcout => \uart_tx_inst.n29\,
            ltout => OPEN,
            carryin => \uart_tx_inst.n1552\,
            carryout => \uart_tx_inst.n1553\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.sub_5_add_2_10_lut_LC_11_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6499\,
            in2 => \N__8376\,
            in3 => \N__5797\,
            lcout => \uart_tx_inst.n28\,
            ltout => OPEN,
            carryin => \bfn_11_3_0_\,
            carryout => \uart_tx_inst.n1554\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.sub_5_add_2_11_lut_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8347\,
            in2 => \N__5794\,
            in3 => \N__5764\,
            lcout => \uart_tx_inst.n27\,
            ltout => OPEN,
            carryin => \uart_tx_inst.n1554\,
            carryout => \uart_tx_inst.n1555\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.sub_5_add_2_12_lut_LC_11_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5761\,
            in2 => \N__8377\,
            in3 => \N__5731\,
            lcout => \uart_tx_inst.n26\,
            ltout => OPEN,
            carryin => \uart_tx_inst.n1555\,
            carryout => \uart_tx_inst.n1556\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.sub_5_add_2_13_lut_LC_11_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8351\,
            in2 => \N__5728\,
            in3 => \N__5698\,
            lcout => \uart_tx_inst.n25\,
            ltout => OPEN,
            carryin => \uart_tx_inst.n1556\,
            carryout => \uart_tx_inst.n1557\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.sub_5_add_2_14_lut_LC_11_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5695\,
            in2 => \N__8378\,
            in3 => \N__5671\,
            lcout => \uart_tx_inst.n24\,
            ltout => OPEN,
            carryin => \uart_tx_inst.n1557\,
            carryout => \uart_tx_inst.n1558\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.sub_5_add_2_15_lut_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8355\,
            in2 => \N__5668\,
            in3 => \N__5635\,
            lcout => \uart_tx_inst.n23\,
            ltout => OPEN,
            carryin => \uart_tx_inst.n1558\,
            carryout => \uart_tx_inst.n1559\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.sub_5_add_2_16_lut_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6070\,
            in2 => \N__8379\,
            in3 => \N__6040\,
            lcout => \uart_tx_inst.n22\,
            ltout => OPEN,
            carryin => \uart_tx_inst.n1559\,
            carryout => \uart_tx_inst.n1560\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.sub_5_add_2_17_lut_LC_11_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8359\,
            in2 => \N__6037\,
            in3 => \N__6004\,
            lcout => \uart_tx_inst.n21\,
            ltout => OPEN,
            carryin => \uart_tx_inst.n1560\,
            carryout => \uart_tx_inst.n1561\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.sub_5_add_2_18_lut_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6001\,
            in2 => \N__8375\,
            in3 => \N__5968\,
            lcout => \uart_tx_inst.n20\,
            ltout => OPEN,
            carryin => \bfn_11_4_0_\,
            carryout => \uart_tx_inst.n1562\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.sub_5_add_2_19_lut_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8342\,
            in2 => \N__5965\,
            in3 => \N__5932\,
            lcout => \uart_tx_inst.n19\,
            ltout => OPEN,
            carryin => \uart_tx_inst.n1562\,
            carryout => \uart_tx_inst.n1563\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.sub_5_add_2_20_lut_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__8343\,
            in1 => \N__5929\,
            in2 => \_gnd_net_\,
            in3 => \N__5905\,
            lcout => \uart_tx_inst.n18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.add_144_2_lut_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7959\,
            in2 => \_gnd_net_\,
            in3 => \N__5881\,
            lcout => \uart_rx_inst.n328\,
            ltout => OPEN,
            carryin => \bfn_11_5_0_\,
            carryout => \uart_rx_inst.n1530\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.add_144_3_lut_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8241\,
            in2 => \N__7881\,
            in3 => \N__5869\,
            lcout => \uart_rx_inst.n327\,
            ltout => OPEN,
            carryin => \uart_rx_inst.n1530\,
            carryout => \uart_rx_inst.n1531\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.add_144_4_lut_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8245\,
            in2 => \N__7785\,
            in3 => \N__5857\,
            lcout => \uart_rx_inst.n326\,
            ltout => OPEN,
            carryin => \uart_rx_inst.n1531\,
            carryout => \uart_rx_inst.n1532\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.add_144_5_lut_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8242\,
            in2 => \N__8858\,
            in3 => \N__6172\,
            lcout => \uart_rx_inst.n325\,
            ltout => OPEN,
            carryin => \uart_rx_inst.n1532\,
            carryout => \uart_rx_inst.n1533\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.add_144_6_lut_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8246\,
            in2 => \N__8770\,
            in3 => \N__6157\,
            lcout => \uart_rx_inst.n324\,
            ltout => OPEN,
            carryin => \uart_rx_inst.n1533\,
            carryout => \uart_rx_inst.n1534\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.add_144_7_lut_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8243\,
            in2 => \N__8669\,
            in3 => \N__6145\,
            lcout => \uart_rx_inst.n323\,
            ltout => OPEN,
            carryin => \uart_rx_inst.n1534\,
            carryout => \uart_rx_inst.n1535\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.add_144_8_lut_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8247\,
            in2 => \N__8566\,
            in3 => \N__6130\,
            lcout => \uart_rx_inst.n322\,
            ltout => OPEN,
            carryin => \uart_rx_inst.n1535\,
            carryout => \uart_rx_inst.n1536\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.add_144_9_lut_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8244\,
            in2 => \N__8463\,
            in3 => \N__6118\,
            lcout => \uart_rx_inst.n321\,
            ltout => OPEN,
            carryin => \uart_rx_inst.n1536\,
            carryout => \uart_rx_inst.n1537\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.add_144_10_lut_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8262\,
            in2 => \N__7972\,
            in3 => \N__6103\,
            lcout => \uart_rx_inst.n320\,
            ltout => OPEN,
            carryin => \bfn_11_6_0_\,
            carryout => \uart_rx_inst.n1538\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.add_144_11_lut_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8328\,
            in2 => \N__7882\,
            in3 => \N__6088\,
            lcout => \uart_rx_inst.n319\,
            ltout => OPEN,
            carryin => \uart_rx_inst.n1538\,
            carryout => \uart_rx_inst.n1539\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.add_144_12_lut_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8263\,
            in2 => \N__7787\,
            in3 => \N__6073\,
            lcout => \uart_rx_inst.n318\,
            ltout => OPEN,
            carryin => \uart_rx_inst.n1539\,
            carryout => \uart_rx_inst.n1540\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.add_144_13_lut_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8329\,
            in2 => \N__8848\,
            in3 => \N__6400\,
            lcout => \uart_rx_inst.n317\,
            ltout => OPEN,
            carryin => \uart_rx_inst.n1540\,
            carryout => \uart_rx_inst.n1541\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.add_144_14_lut_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8264\,
            in2 => \N__8757\,
            in3 => \N__6385\,
            lcout => \uart_rx_inst.n316\,
            ltout => OPEN,
            carryin => \uart_rx_inst.n1541\,
            carryout => \uart_rx_inst.n1542\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.add_144_15_lut_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8330\,
            in2 => \N__8663\,
            in3 => \N__6370\,
            lcout => \uart_rx_inst.n315\,
            ltout => OPEN,
            carryin => \uart_rx_inst.n1542\,
            carryout => \uart_rx_inst.n1543\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.add_144_16_lut_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8265\,
            in2 => \N__8564\,
            in3 => \N__6355\,
            lcout => \uart_rx_inst.n314\,
            ltout => OPEN,
            carryin => \uart_rx_inst.n1543\,
            carryout => \uart_rx_inst.n1544\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.add_144_17_lut_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8331\,
            in2 => \N__8453\,
            in3 => \N__6340\,
            lcout => \uart_rx_inst.n313\,
            ltout => OPEN,
            carryin => \uart_rx_inst.n1544\,
            carryout => \uart_rx_inst.n1545\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.add_144_18_lut_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8169\,
            in2 => \_gnd_net_\,
            in3 => \N__6337\,
            lcout => \uart_rx_inst.n312\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_inst.i1573_2_lut_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7809\,
            in2 => \_gnd_net_\,
            in3 => \N__6314\,
            lcout => \uart_rx_inst.n1746\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.i13_4_lut_LC_12_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__6873\,
            in1 => \N__6207\,
            in2 => \N__6498\,
            in3 => \N__6849\,
            lcout => \uart_tx_inst.n32_adj_197\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.i737_3_lut_LC_12_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6187\,
            in2 => \N__6832\,
            in3 => \N__6930\,
            lcout => OPEN,
            ltout => \uart_tx_inst.n865_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.prescale_reg__i4_LC_12_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__7877\,
            in1 => \N__6597\,
            in2 => \N__6880\,
            in3 => \N__6725\,
            lcout => \uart_tx_inst.prescale_reg_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7384\,
            ce => \N__6475\,
            sr => \N__7227\
        );

    \uart_tx_inst.i742_3_lut_LC_12_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6811\,
            in2 => \N__6862\,
            in3 => \N__6897\,
            lcout => OPEN,
            ltout => \uart_tx_inst.n870_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.prescale_reg__i5_LC_12_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__6726\,
            in1 => \N__7788\,
            in2 => \N__6853\,
            in3 => \N__6603\,
            lcout => \uart_tx_inst.prescale_reg_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7384\,
            ce => \N__6475\,
            sr => \N__7227\
        );

    \uart_tx_inst.i757_3_lut_LC_12_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__8055\,
            in1 => \N__6812\,
            in2 => \_gnd_net_\,
            in3 => \N__6736\,
            lcout => OPEN,
            ltout => \uart_tx_inst.n885_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.prescale_reg__i8_LC_12_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__6727\,
            in1 => \N__8667\,
            in2 => \N__6607\,
            in3 => \N__6604\,
            lcout => \uart_tx_inst.prescale_reg_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7384\,
            ce => \N__6475\,
            sr => \N__7227\
        );

    \uart_tx_inst.data_reg_i0_i0_LC_12_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__7650\,
            in1 => \N__6424\,
            in2 => \N__7939\,
            in3 => \N__7520\,
            lcout => \uart_tx_inst.data_reg_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7383\,
            ce => \N__7546\,
            sr => \_gnd_net_\
        );

    \uart_tx_inst.data_reg_i0_i1_LC_12_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__7521\,
            in1 => \N__7651\,
            in2 => \N__7884\,
            in3 => \N__6418\,
            lcout => \uart_tx_inst.data_reg_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7383\,
            ce => \N__7546\,
            sr => \_gnd_net_\
        );

    \uart_tx_inst.data_reg_i0_i2_LC_12_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__7652\,
            in1 => \N__7687\,
            in2 => \N__7789\,
            in3 => \N__7522\,
            lcout => \uart_tx_inst.data_reg_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7383\,
            ce => \N__7546\,
            sr => \_gnd_net_\
        );

    \uart_tx_inst.data_reg_i0_i3_LC_12_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__7523\,
            in1 => \N__7653\,
            in2 => \N__8867\,
            in3 => \N__7681\,
            lcout => \uart_tx_inst.data_reg_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7383\,
            ce => \N__7546\,
            sr => \_gnd_net_\
        );

    \uart_tx_inst.data_reg_i0_i4_LC_12_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__7654\,
            in1 => \N__8771\,
            in2 => \N__7675\,
            in3 => \N__7524\,
            lcout => \uart_tx_inst.data_reg_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7383\,
            ce => \N__7546\,
            sr => \_gnd_net_\
        );

    \uart_tx_inst.data_reg_i0_i5_LC_12_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__7525\,
            in1 => \N__7655\,
            in2 => \N__8673\,
            in3 => \N__7666\,
            lcout => \uart_tx_inst.data_reg_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7383\,
            ce => \N__7546\,
            sr => \_gnd_net_\
        );

    \uart_tx_inst.data_reg_i0_i6_LC_12_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__7656\,
            in1 => \N__7552\,
            in2 => \N__8572\,
            in3 => \N__7526\,
            lcout => \uart_tx_inst.data_reg_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7383\,
            ce => \N__7546\,
            sr => \_gnd_net_\
        );

    \uart_tx_inst.data_reg_i0_i7_LC_12_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__7527\,
            in1 => \N__7657\,
            in2 => \N__8458\,
            in3 => \N__7570\,
            lcout => \uart_tx_inst.data_reg_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7383\,
            ce => \N__7546\,
            sr => \_gnd_net_\
        );

    \uart_tx_inst.txd_reg_50_LC_12_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__7534\,
            in1 => \N__7528\,
            in2 => \_gnd_net_\,
            in3 => \N__7441\,
            lcout => txd_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7381\,
            ce => \N__7279\,
            sr => \N__7262\
        );

    \uart_tx_inst.sub_8_add_2_2_lut_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7958\,
            in2 => \_gnd_net_\,
            in3 => \N__6937\,
            lcout => n108,
            ltout => OPEN,
            carryin => \bfn_12_5_0_\,
            carryout => \uart_tx_inst.n1582\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.sub_8_add_2_3_lut_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8255\,
            in2 => \N__7846\,
            in3 => \N__6907\,
            lcout => n107,
            ltout => OPEN,
            carryin => \uart_tx_inst.n1582\,
            carryout => \uart_tx_inst.n1583\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.sub_8_add_2_4_lut_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8259\,
            in2 => \N__7750\,
            in3 => \N__8110\,
            lcout => n106,
            ltout => OPEN,
            carryin => \uart_tx_inst.n1583\,
            carryout => \uart_tx_inst.n1584\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.sub_8_add_2_5_lut_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8256\,
            in2 => \N__8847\,
            in3 => \N__8083\,
            lcout => n105,
            ltout => OPEN,
            carryin => \uart_tx_inst.n1584\,
            carryout => \uart_tx_inst.n1585\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.sub_8_add_2_6_lut_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8260\,
            in2 => \N__8753\,
            in3 => \N__8059\,
            lcout => n104,
            ltout => OPEN,
            carryin => \uart_tx_inst.n1585\,
            carryout => \uart_tx_inst.n1586\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.sub_8_add_2_7_lut_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8257\,
            in2 => \N__8668\,
            in3 => \N__8032\,
            lcout => n103,
            ltout => OPEN,
            carryin => \uart_tx_inst.n1586\,
            carryout => \uart_tx_inst.n1587\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.sub_8_add_2_8_lut_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8261\,
            in2 => \N__8565\,
            in3 => \N__8005\,
            lcout => n102,
            ltout => OPEN,
            carryin => \uart_tx_inst.n1587\,
            carryout => \uart_tx_inst.n1588\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.sub_8_add_2_9_lut_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8258\,
            in2 => \N__8454\,
            in3 => \N__7975\,
            lcout => n101,
            ltout => OPEN,
            carryin => \uart_tx_inst.n1588\,
            carryout => \uart_tx_inst.n1589\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.sub_8_add_2_10_lut_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8332\,
            in2 => \N__7971\,
            in3 => \N__7888\,
            lcout => n100,
            ltout => OPEN,
            carryin => \bfn_12_6_0_\,
            carryout => \uart_tx_inst.n1590\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.sub_8_add_2_11_lut_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8266\,
            in2 => \N__7885\,
            in3 => \N__7792\,
            lcout => n99,
            ltout => OPEN,
            carryin => \uart_tx_inst.n1590\,
            carryout => \uart_tx_inst.n1591\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.sub_8_add_2_12_lut_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8333\,
            in2 => \N__7786\,
            in3 => \N__7690\,
            lcout => n98,
            ltout => OPEN,
            carryin => \uart_tx_inst.n1591\,
            carryout => \uart_tx_inst.n1592\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.sub_8_add_2_13_lut_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8267\,
            in2 => \N__8835\,
            in3 => \N__8779\,
            lcout => n97,
            ltout => OPEN,
            carryin => \uart_tx_inst.n1592\,
            carryout => \uart_tx_inst.n1593\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.sub_8_add_2_14_lut_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8334\,
            in2 => \N__8741\,
            in3 => \N__8677\,
            lcout => n96,
            ltout => OPEN,
            carryin => \uart_tx_inst.n1593\,
            carryout => \uart_tx_inst.n1594\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.sub_8_add_2_15_lut_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8268\,
            in2 => \N__8626\,
            in3 => \N__8575\,
            lcout => n95,
            ltout => OPEN,
            carryin => \uart_tx_inst.n1594\,
            carryout => \uart_tx_inst.n1595\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.sub_8_add_2_16_lut_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8335\,
            in2 => \N__8528\,
            in3 => \N__8467\,
            lcout => n94,
            ltout => OPEN,
            carryin => \uart_tx_inst.n1595\,
            carryout => \uart_tx_inst.n1596\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx_inst.sub_8_add_2_17_lut_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__8434\,
            in1 => \N__8269\,
            in2 => \_gnd_net_\,
            in3 => \N__8134\,
            lcout => n93,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
